-- Version: v11.8 11.8.0.26

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreAPB3 is

    port( m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(15 downto 12);
          CoreAPB3_0_APBmslave0_PSELx            : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx : in    std_logic
        );

end CoreAPB3;

architecture DEF_ARCH of CoreAPB3 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \iPSELS_raw_1[0]_net_1\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \iPSELS_raw_1[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15), B
         => m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14), Y => 
        \iPSELS_raw_1[0]_net_1\);
    
    \iPSELS_raw[0]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx, B => 
        \iPSELS_raw_1[0]_net_1\, C => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13), D => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12), Y => 
        CoreAPB3_0_APBmslave0_PSELx);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_CommsFPGA_CCC_0_FCCC is

    port( m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : in    std_logic;
          CommsFPGA_CCC_0_LOCK                      : out   std_logic;
          CommsFPGA_CCC_0_GL1                       : out   std_logic;
          CommsFPGA_CCC_0_GL0                       : out   std_logic
        );

end m2s010_som_CommsFPGA_CCC_0_FCCC;

architecture DEF_ARCH of m2s010_som_CommsFPGA_CCC_0_FCCC is 

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CCC

            generic (INIT:std_logic_vector(209 downto 0) := "00" & x"0000000000000000000000000000000000000000000000000000"; 
        VCOFREQUENCY:real := 0.0);

    port( Y0              : out   std_logic;
          Y1              : out   std_logic;
          Y2              : out   std_logic;
          Y3              : out   std_logic;
          PRDATA          : out   std_logic_vector(7 downto 0);
          LOCK            : out   std_logic;
          BUSY            : out   std_logic;
          CLK0            : in    std_logic := 'U';
          CLK1            : in    std_logic := 'U';
          CLK2            : in    std_logic := 'U';
          CLK3            : in    std_logic := 'U';
          NGMUX0_SEL      : in    std_logic := 'U';
          NGMUX1_SEL      : in    std_logic := 'U';
          NGMUX2_SEL      : in    std_logic := 'U';
          NGMUX3_SEL      : in    std_logic := 'U';
          NGMUX0_HOLD_N   : in    std_logic := 'U';
          NGMUX1_HOLD_N   : in    std_logic := 'U';
          NGMUX2_HOLD_N   : in    std_logic := 'U';
          NGMUX3_HOLD_N   : in    std_logic := 'U';
          NGMUX0_ARST_N   : in    std_logic := 'U';
          NGMUX1_ARST_N   : in    std_logic := 'U';
          NGMUX2_ARST_N   : in    std_logic := 'U';
          NGMUX3_ARST_N   : in    std_logic := 'U';
          PLL_BYPASS_N    : in    std_logic := 'U';
          PLL_ARST_N      : in    std_logic := 'U';
          PLL_POWERDOWN_N : in    std_logic := 'U';
          GPD0_ARST_N     : in    std_logic := 'U';
          GPD1_ARST_N     : in    std_logic := 'U';
          GPD2_ARST_N     : in    std_logic := 'U';
          GPD3_ARST_N     : in    std_logic := 'U';
          PRESET_N        : in    std_logic := 'U';
          PCLK            : in    std_logic := 'U';
          PSEL            : in    std_logic := 'U';
          PENABLE         : in    std_logic := 'U';
          PWRITE          : in    std_logic := 'U';
          PADDR           : in    std_logic_vector(7 downto 2) := (others => 'U');
          PWDATA          : in    std_logic_vector(7 downto 0) := (others => 'U');
          CLK0_PAD        : in    std_logic := 'U';
          CLK1_PAD        : in    std_logic := 'U';
          CLK2_PAD        : in    std_logic := 'U';
          CLK3_PAD        : in    std_logic := 'U';
          GL0             : out   std_logic;
          GL1             : out   std_logic;
          GL2             : out   std_logic;
          GL3             : out   std_logic;
          RCOSC_25_50MHZ  : in    std_logic := 'U';
          RCOSC_1MHZ      : in    std_logic := 'U';
          XTLOSC          : in    std_logic := 'U'
        );
  end component;

    signal GL0_net, GL1_net, VCC_net_1, GND_net_1 : std_logic;
    signal nc8, nc7, nc6, nc2, nc5, nc4, nc3, nc1 : std_logic;

begin 


    GL1_INST : CLKINT
      port map(A => GL1_net, Y => CommsFPGA_CCC_0_GL1);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    GL0_INST : CLKINT
      port map(A => GL0_net, Y => CommsFPGA_CCC_0_GL0);
    
    CCC_INST : CCC

              generic map(INIT => "00" & x"000007FB8000044164000F18C6309C231839DE40404C41803000",
         VCOFREQUENCY => 980.0)

      port map(Y0 => OPEN, Y1 => OPEN, Y2 => OPEN, Y3 => OPEN, 
        PRDATA(7) => nc8, PRDATA(6) => nc7, PRDATA(5) => nc6, 
        PRDATA(4) => nc2, PRDATA(3) => nc5, PRDATA(2) => nc4, 
        PRDATA(1) => nc3, PRDATA(0) => nc1, LOCK => 
        CommsFPGA_CCC_0_LOCK, BUSY => OPEN, CLK0 => VCC_net_1, 
        CLK1 => VCC_net_1, CLK2 => VCC_net_1, CLK3 => VCC_net_1, 
        NGMUX0_SEL => GND_net_1, NGMUX1_SEL => GND_net_1, 
        NGMUX2_SEL => GND_net_1, NGMUX3_SEL => GND_net_1, 
        NGMUX0_HOLD_N => VCC_net_1, NGMUX1_HOLD_N => VCC_net_1, 
        NGMUX2_HOLD_N => VCC_net_1, NGMUX3_HOLD_N => VCC_net_1, 
        NGMUX0_ARST_N => VCC_net_1, NGMUX1_ARST_N => VCC_net_1, 
        NGMUX2_ARST_N => VCC_net_1, NGMUX3_ARST_N => VCC_net_1, 
        PLL_BYPASS_N => VCC_net_1, PLL_ARST_N => VCC_net_1, 
        PLL_POWERDOWN_N => VCC_net_1, GPD0_ARST_N => VCC_net_1, 
        GPD1_ARST_N => VCC_net_1, GPD2_ARST_N => VCC_net_1, 
        GPD3_ARST_N => VCC_net_1, PRESET_N => GND_net_1, PCLK => 
        VCC_net_1, PSEL => VCC_net_1, PENABLE => VCC_net_1, 
        PWRITE => VCC_net_1, PADDR(7) => VCC_net_1, PADDR(6) => 
        VCC_net_1, PADDR(5) => VCC_net_1, PADDR(4) => VCC_net_1, 
        PADDR(3) => VCC_net_1, PADDR(2) => VCC_net_1, PWDATA(7)
         => VCC_net_1, PWDATA(6) => VCC_net_1, PWDATA(5) => 
        VCC_net_1, PWDATA(4) => VCC_net_1, PWDATA(3) => VCC_net_1, 
        PWDATA(2) => VCC_net_1, PWDATA(1) => VCC_net_1, PWDATA(0)
         => VCC_net_1, CLK0_PAD => GND_net_1, CLK1_PAD => 
        GND_net_1, CLK2_PAD => GND_net_1, CLK3_PAD => GND_net_1, 
        GL0 => GL0_net, GL1 => GL1_net, GL2 => OPEN, GL3 => OPEN, 
        RCOSC_25_50MHZ => GND_net_1, RCOSC_1MHZ => GND_net_1, 
        XTLOSC => m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_ID_RES_0_IO is

    port( ID_RES  : in    std_logic_vector(3 downto 0);
          Y_net_0 : out   std_logic_vector(3 downto 0)
        );

end m2s010_som_ID_RES_0_IO;

architecture DEF_ARCH of m2s010_som_ID_RES_0_IO is 

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : INBUF
      port map(PAD => ID_RES(0), Y => Y_net_0(0));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    U0_3 : INBUF
      port map(PAD => ID_RES(3), Y => Y_net_0(3));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    U0_2 : INBUF
      port map(PAD => ID_RES(2), Y => Y_net_0(2));
    
    U0_1 : INBUF
      port map(PAD => ID_RES(1), Y => Y_net_0(1));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_GPIO_1_IO is

    port( GPIO_1_BI_0                       : inout std_logic := 'Z';
          GPIO_1_in_0                       : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_1_M2F_OE : in    std_logic;
          GPIO_1_M2F                        : in    std_logic
        );

end m2s010_som_sb_GPIO_1_IO;

architecture DEF_ARCH of m2s010_som_sb_GPIO_1_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      generic map(IOSTD => "LVCMOS33")

      port map(PAD => GPIO_1_BI_0, D => GPIO_1_M2F, E => 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE, Y => GPIO_1_in_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_CAM_SPI_1_CLK_IO is

    port( CAM_SPI_1_CLK_Y_0                    : out   std_logic;
          SPI_1_CLK_0                          : inout std_logic := 'Z';
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic;
          m2s010_som_sb_MSS_0_SPI_1_CLK_M2F    : in    std_logic
        );

end m2s010_som_sb_CAM_SPI_1_CLK_IO;

architecture DEF_ARCH of m2s010_som_sb_CAM_SPI_1_CLK_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      port map(PAD => SPI_1_CLK_0, D => 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F, E => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, Y => 
        CAM_SPI_1_CLK_Y_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_GPIO_7_IO is

    port( GPIO_7_PADI_0                     : inout std_logic := 'Z';
          GPIO_7_Y_0                        : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F_OE : in    std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F    : in    std_logic
        );

end m2s010_som_sb_GPIO_7_IO;

architecture DEF_ARCH of m2s010_som_sb_GPIO_7_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      port map(PAD => GPIO_7_PADI_0, D => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F, E => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE, Y => GPIO_7_Y_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_CAM_SPI_1_SS0_IO is

    port( SPI_1_SS0_CAM_0                      : inout std_logic := 'Z';
          CAM_SPI_1_SS0_Y_0                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F    : in    std_logic
        );

end m2s010_som_sb_CAM_SPI_1_SS0_IO;

architecture DEF_ARCH of m2s010_som_sb_CAM_SPI_1_SS0_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      port map(PAD => SPI_1_SS0_CAM_0, D => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F, E => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, Y => 
        CAM_SPI_1_SS0_Y_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_MSS is

    port( CORECONFIGP_0_MDDR_APBmslave_PWDATA              : in    std_logic_vector(15 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PADDR               : in    std_logic_vector(10 downto 2);
          MAC_MII_RXD_c                                    : in    std_logic_vector(3 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA  : in    std_logic_vector(17 downto 0);
          Y_net_0                                          : in    std_logic_vector(3 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA_m                   : in    std_logic_vector(7 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PRDATA              : out   std_logic_vector(15 downto 0);
          MAC_MII_TXD_c                                    : out   std_logic_vector(3 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA  : out   std_logic_vector(16 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR   : out   std_logic_vector(15 downto 2);
          CoreAPB3_0_APBmslave0_PWDATA                     : out   std_logic_vector(7 downto 0);
          m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR           : out   std_logic_vector(15 downto 12);
          CoreAPB3_0_APBmslave0_PADDR                      : out   std_logic_vector(7 downto 0);
          MDDR_ADDR                                        : out   std_logic_vector(15 downto 0);
          MDDR_BA                                          : out   std_logic_vector(2 downto 0);
          MDDR_DM_RDQS                                     : inout std_logic_vector(1 downto 0) := (others => 'Z');
          MDDR_DQ                                          : inout std_logic_vector(15 downto 0) := (others => 'Z');
          MDDR_DQS                                         : inout std_logic_vector(1 downto 0) := (others => 'Z');
          CAM_SPI_1_CLK_Y_0                                : in    std_logic;
          GPIO_7_Y_0                                       : in    std_logic;
          GPIO_6_Y_0                                       : in    std_logic;
          DEBOUNCE_OUT_net_0_0                             : in    std_logic;
          GPIO_1_in_0                                      : in    std_logic;
          MDDR_CLK                                         : out   std_logic;
          MDDR_CLK_N                                       : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PWRITE              : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PSELx               : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PENABLE             : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz                        : in    std_logic;
          MAC_MII_TX_CLK_c                                 : in    std_logic;
          SPI_1_SS0_MX_Y                                   : in    std_logic;
          SPI_1_DI                                         : in    std_logic;
          MAC_MII_RX_ER_c                                  : in    std_logic;
          MAC_MII_RX_DV_c                                  : in    std_logic;
          MAC_MII_RX_CLK_c                                 : in    std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR : in    std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY  : in    std_logic;
          MMUART_0_RXD_F2M_c                               : in    std_logic;
          DEBOUNCE_OUT_2_c                                 : in    std_logic;
          DEBOUNCE_OUT_1_c                                 : in    std_logic;
          BIBUF_0_Y                                        : in    std_logic;
          FAB_CCC_LOCK                                     : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY_i_m_i               : in    std_logic;
          CommsFPGA_top_0_INT                              : in    std_logic;
          MAC_MII_CRS_c                                    : in    std_logic;
          MAC_MII_COL_c                                    : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PSLVERR             : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PREADY              : out   std_logic;
          MAC_MII_TX_EN_c                                  : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE             : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F                : out   std_logic;
          SPI_1_DO_CAM_c                                   : out   std_logic;
          GPIO_11_M2F_c                                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_CLK_M2F                : out   std_logic;
          GPIO_8_M2F_c                                     : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F                   : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F_OE                : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F                   : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F_OE                : out   std_logic;
          GPIO_5_M2F_c                                     : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE  : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx   : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE : out   std_logic;
          GPIO_24_M2F_c                                    : out   std_logic;
          MMUART_0_TXD_M2F_c                               : out   std_logic;
          m2s010_som_sb_0_GPIO_28_SW_RESET                 : out   std_logic;
          GPIO_21_M2F_c                                    : out   std_logic;
          GPIO_22_M2F_c                                    : out   std_logic;
          m2s010_som_sb_MSS_0_MAC_MII_MDO                  : out   std_logic;
          m2s010_som_sb_MSS_0_MAC_MII_MDO_EN               : out   std_logic;
          MAC_MII_MDC_c                                    : out   std_logic;
          GPIO_1_M2F                                       : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_1_M2F_OE                : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F          : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE                     : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx           : out   std_logic;
          CoreAPB3_0_APBmslave0_PENABLE                    : out   std_logic;
          GPIO_0_BI                                        : inout std_logic := 'Z';
          GPIO_3_BI                                        : inout std_logic := 'Z';
          GPIO_4_BI                                        : inout std_logic := 'Z';
          GPIO_12_BI                                       : inout std_logic := 'Z';
          GPIO_14_BI                                       : inout std_logic := 'Z';
          GPIO_15_BI                                       : inout std_logic := 'Z';
          GPIO_16_BI                                       : inout std_logic := 'Z';
          GPIO_17_BI                                       : inout std_logic := 'Z';
          GPIO_18_BI                                       : inout std_logic := 'Z';
          GPIO_20_OUT                                      : out   std_logic;
          GPIO_25_BI                                       : inout std_logic := 'Z';
          GPIO_26_BI                                       : inout std_logic := 'Z';
          GPIO_31_BI                                       : inout std_logic := 'Z';
          I2C_1_SCL                                        : inout std_logic := 'Z';
          I2C_1_SDA                                        : inout std_logic := 'Z';
          MDDR_CAS_N                                       : out   std_logic;
          MDDR_CKE                                         : out   std_logic;
          MDDR_CS_N                                        : out   std_logic;
          MDDR_DQS_TMATCH_0_IN                             : in    std_logic;
          MDDR_DQS_TMATCH_0_OUT                            : out   std_logic;
          MDDR_ODT                                         : out   std_logic;
          MDDR_RAS_N                                       : out   std_logic;
          MDDR_RESET_N                                     : out   std_logic;
          MDDR_WE_N                                        : out   std_logic;
          MMUART_1_RXD                                     : in    std_logic;
          MMUART_1_TXD                                     : out   std_logic;
          SPI_0_CLK                                        : inout std_logic := 'Z';
          SPI_0_DI                                         : in    std_logic;
          SPI_0_DO                                         : out   std_logic;
          SPI_0_SS0                                        : inout std_logic := 'Z';
          SPI_0_SS1                                        : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK_i                       : out   std_logic;
          CORECONFIGP_0_APB_S_PRESET_N                     : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK                         : out   std_logic
        );

end m2s010_som_sb_MSS;

architecture DEF_ARCH of m2s010_som_sb_MSS is 

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component TRIBUFF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component MSS_060

            generic (INIT:std_logic_vector(1437 downto 0) := "00" & x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"; 
        ACT_UBITS:std_logic_vector(55 downto 0) := x"FFFFFFFFFFFFFF"; 
        MEMORYFILE:string := ""; RTC_MAIN_XTL_FREQ:real := 0.0; 
        RTC_MAIN_XTL_MODE:string := "1"; DDR_CLK_FREQ:real := 0.0
        );

    port( CAN_RXBUS_MGPIO3A_H2F_A                 : out   std_logic;
          CAN_RXBUS_MGPIO3A_H2F_B                 : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_A                : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_B                : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_A                 : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_B                 : out   std_logic;
          CLK_CONFIG_APB                          : out   std_logic;
          COMMS_INT                               : out   std_logic;
          CONFIG_PRESET_N                         : out   std_logic;
          EDAC_ERROR                              : out   std_logic_vector(7 downto 0);
          F_FM0_RDATA                             : out   std_logic_vector(31 downto 0);
          F_FM0_READYOUT                          : out   std_logic;
          F_FM0_RESP                              : out   std_logic;
          F_HM0_ADDR                              : out   std_logic_vector(31 downto 0);
          F_HM0_ENABLE                            : out   std_logic;
          F_HM0_SEL                               : out   std_logic;
          F_HM0_SIZE                              : out   std_logic_vector(1 downto 0);
          F_HM0_TRANS1                            : out   std_logic;
          F_HM0_WDATA                             : out   std_logic_vector(31 downto 0);
          F_HM0_WRITE                             : out   std_logic;
          FAB_CHRGVBUS                            : out   std_logic;
          FAB_DISCHRGVBUS                         : out   std_logic;
          FAB_DMPULLDOWN                          : out   std_logic;
          FAB_DPPULLDOWN                          : out   std_logic;
          FAB_DRVVBUS                             : out   std_logic;
          FAB_IDPULLUP                            : out   std_logic;
          FAB_OPMODE                              : out   std_logic_vector(1 downto 0);
          FAB_SUSPENDM                            : out   std_logic;
          FAB_TERMSEL                             : out   std_logic;
          FAB_TXVALID                             : out   std_logic;
          FAB_VCONTROL                            : out   std_logic_vector(3 downto 0);
          FAB_VCONTROLLOADM                       : out   std_logic;
          FAB_XCVRSEL                             : out   std_logic_vector(1 downto 0);
          FAB_XDATAOUT                            : out   std_logic_vector(7 downto 0);
          FACC_GLMUX_SEL                          : out   std_logic;
          FIC32_0_MASTER                          : out   std_logic_vector(1 downto 0);
          FIC32_1_MASTER                          : out   std_logic_vector(1 downto 0);
          FPGA_RESET_N                            : out   std_logic;
          GTX_CLK                                 : out   std_logic;
          H2F_INTERRUPT                           : out   std_logic_vector(15 downto 0);
          H2F_NMI                                 : out   std_logic;
          H2FCALIB                                : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_A                 : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_B                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_A                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_B                 : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_A                  : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_B                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_A                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_B                  : out   std_logic;
          MDCF                                    : out   std_logic;
          MDOENF                                  : out   std_logic;
          MDOF                                    : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_A              : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_B              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_A              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_B              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_A              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_B              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_A              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_B              : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_A               : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_B               : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_A              : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_B              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_A              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_B              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_A              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_B              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_A              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_B              : out   std_logic;
          MMUART1_DTR_MGPIO12B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_B              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_A              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_B              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_A              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_B              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_A              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_B              : out   std_logic;
          MPLL_LOCK                               : out   std_logic;
          PER2_FABRIC_PADDR                       : out   std_logic_vector(15 downto 2);
          PER2_FABRIC_PENABLE                     : out   std_logic;
          PER2_FABRIC_PSEL                        : out   std_logic;
          PER2_FABRIC_PWDATA                      : out   std_logic_vector(31 downto 0);
          PER2_FABRIC_PWRITE                      : out   std_logic;
          RTC_MATCH                               : out   std_logic;
          SLEEPDEEP                               : out   std_logic;
          SLEEPHOLDACK                            : out   std_logic;
          SLEEPING                                : out   std_logic;
          SMBALERT_NO0                            : out   std_logic;
          SMBALERT_NO1                            : out   std_logic;
          SMBSUS_NO0                              : out   std_logic;
          SMBSUS_NO1                              : out   std_logic;
          SPI0_CLK_OUT                            : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_A                  : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_B                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_A                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_B                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_A                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_B                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_A                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_B                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_A                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_B                  : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_A                 : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_B                 : out   std_logic;
          SPI0_SS4_MGPIO19A_H2F_A                 : out   std_logic;
          SPI0_SS5_MGPIO20A_H2F_A                 : out   std_logic;
          SPI0_SS6_MGPIO21A_H2F_A                 : out   std_logic;
          SPI0_SS7_MGPIO22A_H2F_A                 : out   std_logic;
          SPI1_CLK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_A                 : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_B                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_A                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_B                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_A                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_B                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_A                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_B                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_A                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_B                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_A                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_B                 : out   std_logic;
          SPI1_SS4_MGPIO17A_H2F_A                 : out   std_logic;
          SPI1_SS5_MGPIO18A_H2F_A                 : out   std_logic;
          SPI1_SS6_MGPIO23A_H2F_A                 : out   std_logic;
          SPI1_SS7_MGPIO24A_H2F_A                 : out   std_logic;
          TCGF                                    : out   std_logic_vector(9 downto 0);
          TRACECLK                                : out   std_logic;
          TRACEDATA                               : out   std_logic_vector(3 downto 0);
          TX_CLK                                  : out   std_logic;
          TX_ENF                                  : out   std_logic;
          TX_ERRF                                 : out   std_logic;
          TXCTL_EN_RIF                            : out   std_logic;
          TXD_RIF                                 : out   std_logic_vector(3 downto 0);
          TXDF                                    : out   std_logic_vector(7 downto 0);
          TXEV                                    : out   std_logic;
          WDOGTIMEOUT                             : out   std_logic;
          F_ARREADY_HREADYOUT1                    : out   std_logic;
          F_AWREADY_HREADYOUT0                    : out   std_logic;
          F_BID                                   : out   std_logic_vector(3 downto 0);
          F_BRESP_HRESP0                          : out   std_logic_vector(1 downto 0);
          F_BVALID                                : out   std_logic;
          F_RDATA_HRDATA01                        : out   std_logic_vector(63 downto 0);
          F_RID                                   : out   std_logic_vector(3 downto 0);
          F_RLAST                                 : out   std_logic;
          F_RRESP_HRESP1                          : out   std_logic_vector(1 downto 0);
          F_RVALID                                : out   std_logic;
          F_WREADY                                : out   std_logic;
          MDDR_FABRIC_PRDATA                      : out   std_logic_vector(15 downto 0);
          MDDR_FABRIC_PREADY                      : out   std_logic;
          MDDR_FABRIC_PSLVERR                     : out   std_logic;
          CAN_RXBUS_F2H_SCP                       : in    std_logic := 'U';
          CAN_TX_EBL_F2H_SCP                      : in    std_logic := 'U';
          CAN_TXBUS_F2H_SCP                       : in    std_logic := 'U';
          COLF                                    : in    std_logic := 'U';
          CRSF                                    : in    std_logic := 'U';
          F2_DMAREADY                             : in    std_logic_vector(1 downto 0) := (others => 'U');
          F2H_INTERRUPT                           : in    std_logic_vector(15 downto 0) := (others => 'U');
          F2HCALIB                                : in    std_logic := 'U';
          F_DMAREADY                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_ADDR                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_ENABLE                            : in    std_logic := 'U';
          F_FM0_MASTLOCK                          : in    std_logic := 'U';
          F_FM0_READY                             : in    std_logic := 'U';
          F_FM0_SEL                               : in    std_logic := 'U';
          F_FM0_SIZE                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_TRANS1                            : in    std_logic := 'U';
          F_FM0_WDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_WRITE                             : in    std_logic := 'U';
          F_HM0_RDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_HM0_READY                             : in    std_logic := 'U';
          F_HM0_RESP                              : in    std_logic := 'U';
          FAB_AVALID                              : in    std_logic := 'U';
          FAB_HOSTDISCON                          : in    std_logic := 'U';
          FAB_IDDIG                               : in    std_logic := 'U';
          FAB_LINESTATE                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          FAB_M3_RESET_N                          : in    std_logic := 'U';
          FAB_PLL_LOCK                            : in    std_logic := 'U';
          FAB_RXACTIVE                            : in    std_logic := 'U';
          FAB_RXERROR                             : in    std_logic := 'U';
          FAB_RXVALID                             : in    std_logic := 'U';
          FAB_RXVALIDH                            : in    std_logic := 'U';
          FAB_SESSEND                             : in    std_logic := 'U';
          FAB_TXREADY                             : in    std_logic := 'U';
          FAB_VBUSVALID                           : in    std_logic := 'U';
          FAB_VSTATUS                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          FAB_XDATAIN                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          GTX_CLKPF                               : in    std_logic := 'U';
          I2C0_BCLK                               : in    std_logic := 'U';
          I2C0_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C0_SDA_F2H_SCP                        : in    std_logic := 'U';
          I2C1_BCLK                               : in    std_logic := 'U';
          I2C1_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C1_SDA_F2H_SCP                        : in    std_logic := 'U';
          MDIF                                    : in    std_logic := 'U';
          MGPIO0A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO10A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO12A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO13A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO14A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO15A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO16A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO17B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO18B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO19B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO1A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO20B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO21B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO22B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO24B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO25B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO26B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO27B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO28B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO29B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO2A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO30B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO31B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO3A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO4A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO5A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO6A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO7A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO8A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO9A_F2H_GPIN                        : in    std_logic := 'U';
          MMUART0_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DTR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART0_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_TXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART1_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_TXD_F2H_SCP                     : in    std_logic := 'U';
          PER2_FABRIC_PRDATA                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          PER2_FABRIC_PREADY                      : in    std_logic := 'U';
          PER2_FABRIC_PSLVERR                     : in    std_logic := 'U';
          RCGF                                    : in    std_logic_vector(9 downto 0) := (others => 'U');
          RX_CLKPF                                : in    std_logic := 'U';
          RX_DVF                                  : in    std_logic := 'U';
          RX_ERRF                                 : in    std_logic := 'U';
          RX_EV                                   : in    std_logic := 'U';
          RXDF                                    : in    std_logic_vector(7 downto 0) := (others => 'U');
          SLEEPHOLDREQ                            : in    std_logic := 'U';
          SMBALERT_NI0                            : in    std_logic := 'U';
          SMBALERT_NI1                            : in    std_logic := 'U';
          SMBSUS_NI0                              : in    std_logic := 'U';
          SMBSUS_NI1                              : in    std_logic := 'U';
          SPI0_CLK_IN                             : in    std_logic := 'U';
          SPI0_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS3_F2H_SCP                        : in    std_logic := 'U';
          SPI1_CLK_IN                             : in    std_logic := 'U';
          SPI1_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS3_F2H_SCP                        : in    std_logic := 'U';
          TX_CLKPF                                : in    std_logic := 'U';
          USER_MSS_GPIO_RESET_N                   : in    std_logic := 'U';
          USER_MSS_RESET_N                        : in    std_logic := 'U';
          XCLK_FAB                                : in    std_logic := 'U';
          CLK_BASE                                : in    std_logic := 'U';
          CLK_MDDR_APB                            : in    std_logic := 'U';
          F_ARADDR_HADDR1                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_ARBURST_HTRANS1                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARID_HSEL1                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLEN_HBURST1                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLOCK_HMASTLOCK1                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARSIZE_HSIZE1                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARVALID_HWRITE1                       : in    std_logic := 'U';
          F_AWADDR_HADDR0                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_AWBURST_HTRANS0                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWID_HSEL0                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLEN_HBURST0                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLOCK_HMASTLOCK0                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWSIZE_HSIZE0                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWVALID_HWRITE0                       : in    std_logic := 'U';
          F_BREADY                                : in    std_logic := 'U';
          F_RMW_AXI                               : in    std_logic := 'U';
          F_RREADY                                : in    std_logic := 'U';
          F_WDATA_HWDATA01                        : in    std_logic_vector(63 downto 0) := (others => 'U');
          F_WID_HREADY01                          : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_WLAST                                 : in    std_logic := 'U';
          F_WSTRB                                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          F_WVALID                                : in    std_logic := 'U';
          FPGA_MDDR_ARESET_N                      : in    std_logic := 'U';
          MDDR_FABRIC_PADDR                       : in    std_logic_vector(10 downto 2) := (others => 'U');
          MDDR_FABRIC_PENABLE                     : in    std_logic := 'U';
          MDDR_FABRIC_PSEL                        : in    std_logic := 'U';
          MDDR_FABRIC_PWDATA                      : in    std_logic_vector(15 downto 0) := (others => 'U');
          MDDR_FABRIC_PWRITE                      : in    std_logic := 'U';
          PRESET_N                                : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_IN         : in    std_logic := 'U';
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN        : in    std_logic := 'U';
          CAN_TXBUS_USBA_DATA0_MGPIO2A_IN         : in    std_logic := 'U';
          DM_IN                                   : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_DQ_IN                              : in    std_logic_vector(17 downto 0) := (others => 'U');
          DRAM_DQS_IN                             : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_FIFO_WE_IN                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          I2C0_SCL_USBC_DATA1_MGPIO31B_IN         : in    std_logic := 'U';
          I2C0_SDA_USBC_DATA0_MGPIO30B_IN         : in    std_logic := 'U';
          I2C1_SCL_USBA_DATA4_MGPIO1A_IN          : in    std_logic := 'U';
          I2C1_SDA_USBA_DATA3_MGPIO0A_IN          : in    std_logic := 'U';
          MGPIO0B_IN                              : in    std_logic := 'U';
          MGPIO10B_IN                             : in    std_logic := 'U';
          MGPIO1B_IN                              : in    std_logic := 'U';
          MGPIO25A_IN                             : in    std_logic := 'U';
          MGPIO26A_IN                             : in    std_logic := 'U';
          MGPIO27A_IN                             : in    std_logic := 'U';
          MGPIO28A_IN                             : in    std_logic := 'U';
          MGPIO29A_IN                             : in    std_logic := 'U';
          MGPIO2B_IN                              : in    std_logic := 'U';
          MGPIO30A_IN                             : in    std_logic := 'U';
          MGPIO31A_IN                             : in    std_logic := 'U';
          MGPIO3B_IN                              : in    std_logic := 'U';
          MGPIO4B_IN                              : in    std_logic := 'U';
          MGPIO5B_IN                              : in    std_logic := 'U';
          MGPIO6B_IN                              : in    std_logic := 'U';
          MGPIO7B_IN                              : in    std_logic := 'U';
          MGPIO8B_IN                              : in    std_logic := 'U';
          MGPIO9B_IN                              : in    std_logic := 'U';
          MMUART0_CTS_USBC_DATA7_MGPIO19B_IN      : in    std_logic := 'U';
          MMUART0_DCD_MGPIO22B_IN                 : in    std_logic := 'U';
          MMUART0_DSR_MGPIO20B_IN                 : in    std_logic := 'U';
          MMUART0_DTR_USBC_DATA6_MGPIO18B_IN      : in    std_logic := 'U';
          MMUART0_RI_MGPIO21B_IN                  : in    std_logic := 'U';
          MMUART0_RTS_USBC_DATA5_MGPIO17B_IN      : in    std_logic := 'U';
          MMUART0_RXD_USBC_STP_MGPIO28B_IN        : in    std_logic := 'U';
          MMUART0_SCK_USBC_NXT_MGPIO29B_IN        : in    std_logic := 'U';
          MMUART0_TXD_USBC_DIR_MGPIO27B_IN        : in    std_logic := 'U';
          MMUART1_CTS_MGPIO13B_IN                 : in    std_logic := 'U';
          MMUART1_DCD_MGPIO16B_IN                 : in    std_logic := 'U';
          MMUART1_DSR_MGPIO14B_IN                 : in    std_logic := 'U';
          MMUART1_DTR_MGPIO12B_IN                 : in    std_logic := 'U';
          MMUART1_RI_MGPIO15B_IN                  : in    std_logic := 'U';
          MMUART1_RTS_MGPIO11B_IN                 : in    std_logic := 'U';
          MMUART1_RXD_USBC_DATA3_MGPIO26B_IN      : in    std_logic := 'U';
          MMUART1_SCK_USBC_DATA4_MGPIO25B_IN      : in    std_logic := 'U';
          MMUART1_TXD_USBC_DATA2_MGPIO24B_IN      : in    std_logic := 'U';
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN     : in    std_logic := 'U';
          RGMII_MDC_RMII_MDC_IN                   : in    std_logic := 'U';
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN      : in    std_logic := 'U';
          RGMII_RX_CLK_IN                         : in    std_logic := 'U';
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN  : in    std_logic := 'U';
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN      : in    std_logic := 'U';
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN      : in    std_logic := 'U';
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN     : in    std_logic := 'U';
          RGMII_RXD3_USBB_DATA4_IN                : in    std_logic := 'U';
          RGMII_TX_CLK_IN                         : in    std_logic := 'U';
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN     : in    std_logic := 'U';
          RGMII_TXD0_RMII_TXD0_USBB_DIR_IN        : in    std_logic := 'U';
          RGMII_TXD1_RMII_TXD1_USBB_STP_IN        : in    std_logic := 'U';
          RGMII_TXD2_USBB_DATA5_IN                : in    std_logic := 'U';
          RGMII_TXD3_USBB_DATA6_IN                : in    std_logic := 'U';
          SPI0_SCK_USBA_XCLK_IN                   : in    std_logic := 'U';
          SPI0_SDI_USBA_DIR_MGPIO5A_IN            : in    std_logic := 'U';
          SPI0_SDO_USBA_STP_MGPIO6A_IN            : in    std_logic := 'U';
          SPI0_SS0_USBA_NXT_MGPIO7A_IN            : in    std_logic := 'U';
          SPI0_SS1_USBA_DATA5_MGPIO8A_IN          : in    std_logic := 'U';
          SPI0_SS2_USBA_DATA6_MGPIO9A_IN          : in    std_logic := 'U';
          SPI0_SS3_USBA_DATA7_MGPIO10A_IN         : in    std_logic := 'U';
          SPI0_SS4_MGPIO19A_IN                    : in    std_logic := 'U';
          SPI0_SS5_MGPIO20A_IN                    : in    std_logic := 'U';
          SPI0_SS6_MGPIO21A_IN                    : in    std_logic := 'U';
          SPI0_SS7_MGPIO22A_IN                    : in    std_logic := 'U';
          SPI1_SCK_IN                             : in    std_logic := 'U';
          SPI1_SDI_MGPIO11A_IN                    : in    std_logic := 'U';
          SPI1_SDO_MGPIO12A_IN                    : in    std_logic := 'U';
          SPI1_SS0_MGPIO13A_IN                    : in    std_logic := 'U';
          SPI1_SS1_MGPIO14A_IN                    : in    std_logic := 'U';
          SPI1_SS2_MGPIO15A_IN                    : in    std_logic := 'U';
          SPI1_SS3_MGPIO16A_IN                    : in    std_logic := 'U';
          SPI1_SS4_MGPIO17A_IN                    : in    std_logic := 'U';
          SPI1_SS5_MGPIO18A_IN                    : in    std_logic := 'U';
          SPI1_SS6_MGPIO23A_IN                    : in    std_logic := 'U';
          SPI1_SS7_MGPIO24A_IN                    : in    std_logic := 'U';
          USBC_XCLK_IN                            : in    std_logic := 'U';
          USBD_DATA0_IN                           : in    std_logic := 'U';
          USBD_DATA1_IN                           : in    std_logic := 'U';
          USBD_DATA2_IN                           : in    std_logic := 'U';
          USBD_DATA3_IN                           : in    std_logic := 'U';
          USBD_DATA4_IN                           : in    std_logic := 'U';
          USBD_DATA5_IN                           : in    std_logic := 'U';
          USBD_DATA6_IN                           : in    std_logic := 'U';
          USBD_DATA7_MGPIO23B_IN                  : in    std_logic := 'U';
          USBD_DIR_IN                             : in    std_logic := 'U';
          USBD_NXT_IN                             : in    std_logic := 'U';
          USBD_STP_IN                             : in    std_logic := 'U';
          USBD_XCLK_IN                            : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT        : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT       : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT        : out   std_logic;
          DRAM_ADDR                               : out   std_logic_vector(15 downto 0);
          DRAM_BA                                 : out   std_logic_vector(2 downto 0);
          DRAM_CASN                               : out   std_logic;
          DRAM_CKE                                : out   std_logic;
          DRAM_CLK                                : out   std_logic;
          DRAM_CSN                                : out   std_logic;
          DRAM_DM_RDQS_OUT                        : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OUT                             : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OUT                            : out   std_logic_vector(2 downto 0);
          DRAM_FIFO_WE_OUT                        : out   std_logic_vector(1 downto 0);
          DRAM_ODT                                : out   std_logic;
          DRAM_RASN                               : out   std_logic;
          DRAM_RSTN                               : out   std_logic;
          DRAM_WEN                                : out   std_logic;
          I2C0_SCL_USBC_DATA1_MGPIO31B_OUT        : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OUT        : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OUT         : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OUT         : out   std_logic;
          MGPIO0B_OUT                             : out   std_logic;
          MGPIO10B_OUT                            : out   std_logic;
          MGPIO1B_OUT                             : out   std_logic;
          MGPIO25A_OUT                            : out   std_logic;
          MGPIO26A_OUT                            : out   std_logic;
          MGPIO27A_OUT                            : out   std_logic;
          MGPIO28A_OUT                            : out   std_logic;
          MGPIO29A_OUT                            : out   std_logic;
          MGPIO2B_OUT                             : out   std_logic;
          MGPIO30A_OUT                            : out   std_logic;
          MGPIO31A_OUT                            : out   std_logic;
          MGPIO3B_OUT                             : out   std_logic;
          MGPIO4B_OUT                             : out   std_logic;
          MGPIO5B_OUT                             : out   std_logic;
          MGPIO6B_OUT                             : out   std_logic;
          MGPIO7B_OUT                             : out   std_logic;
          MGPIO8B_OUT                             : out   std_logic;
          MGPIO9B_OUT                             : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT     : out   std_logic;
          MMUART0_DCD_MGPIO22B_OUT                : out   std_logic;
          MMUART0_DSR_MGPIO20B_OUT                : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT     : out   std_logic;
          MMUART0_RI_MGPIO21B_OUT                 : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT     : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OUT       : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OUT       : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OUT       : out   std_logic;
          MMUART1_CTS_MGPIO13B_OUT                : out   std_logic;
          MMUART1_DCD_MGPIO16B_OUT                : out   std_logic;
          MMUART1_DSR_MGPIO14B_OUT                : out   std_logic;
          MMUART1_DTR_MGPIO12B_OUT                : out   std_logic;
          MMUART1_RI_MGPIO15B_OUT                 : out   std_logic;
          MMUART1_RTS_MGPIO11B_OUT                : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT     : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT     : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT     : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT    : out   std_logic;
          RGMII_MDC_RMII_MDC_OUT                  : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT     : out   std_logic;
          RGMII_RX_CLK_OUT                        : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT     : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT     : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT    : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OUT               : out   std_logic;
          RGMII_TX_CLK_OUT                        : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT    : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT       : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OUT       : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OUT               : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OUT               : out   std_logic;
          SPI0_SCK_USBA_XCLK_OUT                  : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OUT           : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OUT           : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OUT           : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OUT         : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OUT         : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OUT        : out   std_logic;
          SPI0_SS4_MGPIO19A_OUT                   : out   std_logic;
          SPI0_SS5_MGPIO20A_OUT                   : out   std_logic;
          SPI0_SS6_MGPIO21A_OUT                   : out   std_logic;
          SPI0_SS7_MGPIO22A_OUT                   : out   std_logic;
          SPI1_SCK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_OUT                   : out   std_logic;
          SPI1_SDO_MGPIO12A_OUT                   : out   std_logic;
          SPI1_SS0_MGPIO13A_OUT                   : out   std_logic;
          SPI1_SS1_MGPIO14A_OUT                   : out   std_logic;
          SPI1_SS2_MGPIO15A_OUT                   : out   std_logic;
          SPI1_SS3_MGPIO16A_OUT                   : out   std_logic;
          SPI1_SS4_MGPIO17A_OUT                   : out   std_logic;
          SPI1_SS5_MGPIO18A_OUT                   : out   std_logic;
          SPI1_SS6_MGPIO23A_OUT                   : out   std_logic;
          SPI1_SS7_MGPIO24A_OUT                   : out   std_logic;
          USBC_XCLK_OUT                           : out   std_logic;
          USBD_DATA0_OUT                          : out   std_logic;
          USBD_DATA1_OUT                          : out   std_logic;
          USBD_DATA2_OUT                          : out   std_logic;
          USBD_DATA3_OUT                          : out   std_logic;
          USBD_DATA4_OUT                          : out   std_logic;
          USBD_DATA5_OUT                          : out   std_logic;
          USBD_DATA6_OUT                          : out   std_logic;
          USBD_DATA7_MGPIO23B_OUT                 : out   std_logic;
          USBD_DIR_OUT                            : out   std_logic;
          USBD_NXT_OUT                            : out   std_logic;
          USBD_STP_OUT                            : out   std_logic;
          USBD_XCLK_OUT                           : out   std_logic;
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OE         : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE        : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OE         : out   std_logic;
          DM_OE                                   : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OE                              : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OE                             : out   std_logic_vector(2 downto 0);
          I2C0_SCL_USBC_DATA1_MGPIO31B_OE         : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OE         : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OE          : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OE          : out   std_logic;
          MGPIO0B_OE                              : out   std_logic;
          MGPIO10B_OE                             : out   std_logic;
          MGPIO1B_OE                              : out   std_logic;
          MGPIO25A_OE                             : out   std_logic;
          MGPIO26A_OE                             : out   std_logic;
          MGPIO27A_OE                             : out   std_logic;
          MGPIO28A_OE                             : out   std_logic;
          MGPIO29A_OE                             : out   std_logic;
          MGPIO2B_OE                              : out   std_logic;
          MGPIO30A_OE                             : out   std_logic;
          MGPIO31A_OE                             : out   std_logic;
          MGPIO3B_OE                              : out   std_logic;
          MGPIO4B_OE                              : out   std_logic;
          MGPIO5B_OE                              : out   std_logic;
          MGPIO6B_OE                              : out   std_logic;
          MGPIO7B_OE                              : out   std_logic;
          MGPIO8B_OE                              : out   std_logic;
          MGPIO9B_OE                              : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OE      : out   std_logic;
          MMUART0_DCD_MGPIO22B_OE                 : out   std_logic;
          MMUART0_DSR_MGPIO20B_OE                 : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OE      : out   std_logic;
          MMUART0_RI_MGPIO21B_OE                  : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OE      : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OE        : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OE        : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OE        : out   std_logic;
          MMUART1_CTS_MGPIO13B_OE                 : out   std_logic;
          MMUART1_DCD_MGPIO16B_OE                 : out   std_logic;
          MMUART1_DSR_MGPIO14B_OE                 : out   std_logic;
          MMUART1_DTR_MGPIO12B_OE                 : out   std_logic;
          MMUART1_RI_MGPIO15B_OE                  : out   std_logic;
          MMUART1_RTS_MGPIO11B_OE                 : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OE      : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OE      : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OE      : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE     : out   std_logic;
          RGMII_MDC_RMII_MDC_OE                   : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE      : out   std_logic;
          RGMII_RX_CLK_OE                         : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE  : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE      : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE      : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE     : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OE                : out   std_logic;
          RGMII_TX_CLK_OE                         : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE     : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OE        : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OE        : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OE                : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OE                : out   std_logic;
          SPI0_SCK_USBA_XCLK_OE                   : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OE            : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OE            : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OE            : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OE          : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OE          : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OE         : out   std_logic;
          SPI0_SS4_MGPIO19A_OE                    : out   std_logic;
          SPI0_SS5_MGPIO20A_OE                    : out   std_logic;
          SPI0_SS6_MGPIO21A_OE                    : out   std_logic;
          SPI0_SS7_MGPIO22A_OE                    : out   std_logic;
          SPI1_SCK_OE                             : out   std_logic;
          SPI1_SDI_MGPIO11A_OE                    : out   std_logic;
          SPI1_SDO_MGPIO12A_OE                    : out   std_logic;
          SPI1_SS0_MGPIO13A_OE                    : out   std_logic;
          SPI1_SS1_MGPIO14A_OE                    : out   std_logic;
          SPI1_SS2_MGPIO15A_OE                    : out   std_logic;
          SPI1_SS3_MGPIO16A_OE                    : out   std_logic;
          SPI1_SS4_MGPIO17A_OE                    : out   std_logic;
          SPI1_SS5_MGPIO18A_OE                    : out   std_logic;
          SPI1_SS6_MGPIO23A_OE                    : out   std_logic;
          SPI1_SS7_MGPIO24A_OE                    : out   std_logic;
          USBC_XCLK_OE                            : out   std_logic;
          USBD_DATA0_OE                           : out   std_logic;
          USBD_DATA1_OE                           : out   std_logic;
          USBD_DATA2_OE                           : out   std_logic;
          USBD_DATA3_OE                           : out   std_logic;
          USBD_DATA4_OE                           : out   std_logic;
          USBD_DATA5_OE                           : out   std_logic;
          USBD_DATA6_OE                           : out   std_logic;
          USBD_DATA7_MGPIO23B_OE                  : out   std_logic;
          USBD_DIR_OE                             : out   std_logic;
          USBD_NXT_OE                             : out   std_logic;
          USBD_STP_OE                             : out   std_logic;
          USBD_XCLK_OE                            : out   std_logic
        );
  end component;

  component OUTBUF_DIFF
    generic (IOSTD:string := "");

    port( D    : in    std_logic := 'U';
          PADP : out   std_logic;
          PADN : out   std_logic
        );
  end component;

    signal \CORECONFIGP_0_APB_S_PCLK\, FIC_2_APB_M_PCLK, 
        \CORECONFIGP_0_APB_S_PRESET_N\, CONFIG_PRESET_N, 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OUT, 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OE, 
        SPI_0_SS0_PAD_Y, 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, 
        SPI_0_DI_PAD_Y, SPI_0_CLK_PAD_Y, 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, 
        MMUART_1_RXD_PAD_Y, MSS_ADLIB_INST_DRAM_WEN, 
        MSS_ADLIB_INST_DRAM_RSTN, MSS_ADLIB_INST_DRAM_RASN, 
        MSS_ADLIB_INST_DRAM_ODT, \DRAM_FIFO_WE_OUT_net_0[0]\, 
        MDDR_DQS_TMATCH_0_IN_PAD_Y, MDDR_DQS_1_PAD_Y, 
        \DRAM_DQS_OUT_net_0[1]\, \DRAM_DQS_OE_net_0[1]\, 
        MDDR_DQS_0_PAD_Y, \DRAM_DQS_OUT_net_0[0]\, 
        \DRAM_DQS_OE_net_0[0]\, MDDR_DQ_15_PAD_Y, 
        \DRAM_DQ_OUT_net_0[15]\, \DRAM_DQ_OE_net_0[15]\, 
        MDDR_DQ_14_PAD_Y, \DRAM_DQ_OUT_net_0[14]\, 
        \DRAM_DQ_OE_net_0[14]\, MDDR_DQ_13_PAD_Y, 
        \DRAM_DQ_OUT_net_0[13]\, \DRAM_DQ_OE_net_0[13]\, 
        MDDR_DQ_12_PAD_Y, \DRAM_DQ_OUT_net_0[12]\, 
        \DRAM_DQ_OE_net_0[12]\, MDDR_DQ_11_PAD_Y, 
        \DRAM_DQ_OUT_net_0[11]\, \DRAM_DQ_OE_net_0[11]\, 
        MDDR_DQ_10_PAD_Y, \DRAM_DQ_OUT_net_0[10]\, 
        \DRAM_DQ_OE_net_0[10]\, MDDR_DQ_9_PAD_Y, 
        \DRAM_DQ_OUT_net_0[9]\, \DRAM_DQ_OE_net_0[9]\, 
        MDDR_DQ_8_PAD_Y, \DRAM_DQ_OUT_net_0[8]\, 
        \DRAM_DQ_OE_net_0[8]\, MDDR_DQ_7_PAD_Y, 
        \DRAM_DQ_OUT_net_0[7]\, \DRAM_DQ_OE_net_0[7]\, 
        MDDR_DQ_6_PAD_Y, \DRAM_DQ_OUT_net_0[6]\, 
        \DRAM_DQ_OE_net_0[6]\, MDDR_DQ_5_PAD_Y, 
        \DRAM_DQ_OUT_net_0[5]\, \DRAM_DQ_OE_net_0[5]\, 
        MDDR_DQ_4_PAD_Y, \DRAM_DQ_OUT_net_0[4]\, 
        \DRAM_DQ_OE_net_0[4]\, MDDR_DQ_3_PAD_Y, 
        \DRAM_DQ_OUT_net_0[3]\, \DRAM_DQ_OE_net_0[3]\, 
        MDDR_DQ_2_PAD_Y, \DRAM_DQ_OUT_net_0[2]\, 
        \DRAM_DQ_OE_net_0[2]\, MDDR_DQ_1_PAD_Y, 
        \DRAM_DQ_OUT_net_0[1]\, \DRAM_DQ_OE_net_0[1]\, 
        MDDR_DQ_0_PAD_Y, \DRAM_DQ_OUT_net_0[0]\, 
        \DRAM_DQ_OE_net_0[0]\, MDDR_DM_RDQS_1_PAD_Y, 
        \DRAM_DM_RDQS_OUT_net_0[1]\, \DM_OE_net_0[1]\, 
        MDDR_DM_RDQS_0_PAD_Y, \DRAM_DM_RDQS_OUT_net_0[0]\, 
        \DM_OE_net_0[0]\, MSS_ADLIB_INST_DRAM_CSN, 
        MSS_ADLIB_INST_DRAM_CKE, MSS_ADLIB_INST_DRAM_CASN, 
        \DRAM_BA_net_0[2]\, \DRAM_BA_net_0[1]\, 
        \DRAM_BA_net_0[0]\, \DRAM_ADDR_net_0[15]\, 
        \DRAM_ADDR_net_0[14]\, \DRAM_ADDR_net_0[13]\, 
        \DRAM_ADDR_net_0[12]\, \DRAM_ADDR_net_0[11]\, 
        \DRAM_ADDR_net_0[10]\, \DRAM_ADDR_net_0[9]\, 
        \DRAM_ADDR_net_0[8]\, \DRAM_ADDR_net_0[7]\, 
        \DRAM_ADDR_net_0[6]\, \DRAM_ADDR_net_0[5]\, 
        \DRAM_ADDR_net_0[4]\, \DRAM_ADDR_net_0[3]\, 
        \DRAM_ADDR_net_0[2]\, \DRAM_ADDR_net_0[1]\, 
        \DRAM_ADDR_net_0[0]\, I2C_1_SDA_PAD_Y, 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT, 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE, 
        I2C_1_SCL_PAD_Y, 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT, 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE, 
        GPIO_GPIO_31_BI_PAD_Y, MSS_ADLIB_INST_MGPIO31A_OUT, 
        MSS_ADLIB_INST_MGPIO31A_OE, GPIO_GPIO_26_BI_PAD_Y, 
        MSS_ADLIB_INST_MGPIO26A_OUT, MSS_ADLIB_INST_MGPIO26A_OE, 
        GPIO_GPIO_25_BI_PAD_Y, MSS_ADLIB_INST_MGPIO25A_OUT, 
        MSS_ADLIB_INST_MGPIO25A_OE, 
        MSS_ADLIB_INST_SPI0_SS5_MGPIO20A_OUT, 
        GPIO_GPIO_18_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OUT, 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OE, 
        GPIO_GPIO_17_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OUT, 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OE, 
        GPIO_GPIO_16_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OUT, 
        MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OE, 
        GPIO_GPIO_15_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OUT, 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OE, 
        GPIO_GPIO_14_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OUT, 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OE, 
        GPIO_GPIO_12_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OUT, 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OE, 
        GPIO_GPIO_4_BI_PAD_Y, 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT, 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE, 
        GPIO_GPIO_3_BI_PAD_Y, 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT, 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OE, 
        GPIO_GPIO_0_BI_PAD_Y, MSS_ADLIB_INST_MGPIO0B_OUT, 
        MSS_ADLIB_INST_MGPIO0B_OE, VCC_net_1, GND_net_1, 
        MSS_ADLIB_INST_DRAM_CLK : std_logic;
    signal nc228, nc203, nc216, nc194, nc151, nc23, nc175, nc58, 
        nc116, nc74, nc133, nc238, nc167, nc84, nc39, nc72, nc212, 
        nc205, nc82, nc145, nc181, nc160, nc57, nc156, nc125, 
        nc211, nc73, nc107, nc66, nc83, nc9, nc171, nc54, nc135, 
        nc41, nc100, nc52, nc186, nc29, nc118, nc60, nc141, nc193, 
        nc214, nc240, nc45, nc53, nc121, nc176, nc220, nc158, 
        nc209, nc246, nc162, nc11, nc131, nc96, nc79, nc226, 
        nc146, nc230, nc89, nc119, nc48, nc213, nc126, nc195, 
        nc188, nc242, nc15, nc236, nc102, nc3, nc207, nc47, nc90, 
        nc222, nc159, nc136, nc241, nc178, nc215, nc59, nc221, 
        nc232, nc18, nc44, nc117, nc189, nc164, nc148, nc42, 
        nc231, nc191, nc17, nc2, nc110, nc128, nc244, nc43, nc179, 
        nc157, nc36, nc224, nc61, nc104, nc138, nc14, nc150, 
        nc196, nc234, nc149, nc12, nc219, nc30, nc243, nc187, 
        nc65, nc7, nc129, nc8, nc223, nc13, nc180, nc26, nc177, 
        nc139, nc245, nc233, nc163, nc112, nc68, nc49, nc217, 
        nc170, nc91, nc225, nc5, nc20, nc198, nc147, nc67, nc152, 
        nc127, nc103, nc235, nc76, nc208, nc140, nc86, nc95, 
        nc120, nc165, nc137, nc64, nc19, nc70, nc182, nc62, nc199, 
        nc80, nc130, nc98, nc114, nc56, nc105, nc63, nc172, nc229, 
        nc97, nc161, nc31, nc154, nc50, nc239, nc142, nc94, nc197, 
        nc122, nc35, nc4, nc227, nc92, nc101, nc184, nc200, nc190, 
        nc166, nc132, nc21, nc237, nc93, nc69, nc206, nc174, nc38, 
        nc113, nc218, nc106, nc25, nc1, nc37, nc202, nc144, nc153, 
        nc46, nc71, nc124, nc81, nc201, nc168, nc34, nc28, nc115, 
        nc192, nc134, nc32, nc40, nc99, nc75, nc183, nc85, nc27, 
        nc108, nc16, nc155, nc51, nc33, nc204, nc173, nc169, nc78, 
        nc24, nc88, nc111, nc55, nc10, nc22, nc210, nc185, nc143, 
        nc77, nc6, nc109, nc87, nc123 : std_logic;

begin 

    CORECONFIGP_0_APB_S_PRESET_N <= 
        \CORECONFIGP_0_APB_S_PRESET_N\;
    CORECONFIGP_0_APB_S_PCLK <= \CORECONFIGP_0_APB_S_PCLK\;

    MDDR_ADDR_6_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[6]\, PAD => MDDR_ADDR(6));
    
    MDDR_CAS_N_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_CASN, PAD => MDDR_CAS_N);
    
    MDDR_RESET_N_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_RSTN, PAD => MDDR_RESET_N);
    
    MDDR_ODT_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_ODT, PAD => MDDR_ODT);
    
    GPIO_GPIO_31_BI_PAD : BIBUF
      port map(PAD => GPIO_31_BI, D => 
        MSS_ADLIB_INST_MGPIO31A_OUT, E => 
        MSS_ADLIB_INST_MGPIO31A_OE, Y => GPIO_GPIO_31_BI_PAD_Y);
    
    MDDR_ADDR_11_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[11]\, PAD => MDDR_ADDR(11));
    
    MMUART_1_TXD_PAD : TRIBUFF
      port map(D => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, PAD
         => MMUART_1_TXD);
    
    MDDR_DQ_10_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(10), D => \DRAM_DQ_OUT_net_0[10]\, 
        E => \DRAM_DQ_OE_net_0[10]\, Y => MDDR_DQ_10_PAD_Y);
    
    MDDR_DQ_1_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(1), D => \DRAM_DQ_OUT_net_0[1]\, E
         => \DRAM_DQ_OE_net_0[1]\, Y => MDDR_DQ_1_PAD_Y);
    
    MDDR_ADDR_7_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[7]\, PAD => MDDR_ADDR(7));
    
    MDDR_DQ_11_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(11), D => \DRAM_DQ_OUT_net_0[11]\, 
        E => \DRAM_DQ_OE_net_0[11]\, Y => MDDR_DQ_11_PAD_Y);
    
    MDDR_DQ_9_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(9), D => \DRAM_DQ_OUT_net_0[9]\, E
         => \DRAM_DQ_OE_net_0[9]\, Y => MDDR_DQ_9_PAD_Y);
    
    MSS_ADLIB_INST_RNI1CJ7 : CLKINT
      port map(A => CONFIG_PRESET_N, Y => 
        \CORECONFIGP_0_APB_S_PRESET_N\);
    
    MDDR_DQ_3_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(3), D => \DRAM_DQ_OUT_net_0[3]\, E
         => \DRAM_DQ_OE_net_0[3]\, Y => MDDR_DQ_3_PAD_Y);
    
    GPIO_GPIO_25_BI_PAD : BIBUF
      port map(PAD => GPIO_25_BI, D => 
        MSS_ADLIB_INST_MGPIO25A_OUT, E => 
        MSS_ADLIB_INST_MGPIO25A_OE, Y => GPIO_GPIO_25_BI_PAD_Y);
    
    MDDR_DQ_0_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(0), D => \DRAM_DQ_OUT_net_0[0]\, E
         => \DRAM_DQ_OE_net_0[0]\, Y => MDDR_DQ_0_PAD_Y);
    
    MDDR_ADDR_12_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[12]\, PAD => MDDR_ADDR(12));
    
    GPIO_GPIO_17_BI_PAD : BIBUF
      port map(PAD => GPIO_17_BI, D => 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OUT, E => 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OE, Y => 
        GPIO_GPIO_17_BI_PAD_Y);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    MDDR_DQ_2_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(2), D => \DRAM_DQ_OUT_net_0[2]\, E
         => \DRAM_DQ_OE_net_0[2]\, Y => MDDR_DQ_2_PAD_Y);
    
    MDDR_DQ_12_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(12), D => \DRAM_DQ_OUT_net_0[12]\, 
        E => \DRAM_DQ_OE_net_0[12]\, Y => MDDR_DQ_12_PAD_Y);
    
    MDDR_CKE_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_CKE, PAD => MDDR_CKE);
    
    MDDR_ADDR_2_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[2]\, PAD => MDDR_ADDR(2));
    
    GPIO_GPIO_0_BI_PAD : BIBUF
      port map(PAD => GPIO_0_BI, D => MSS_ADLIB_INST_MGPIO0B_OUT, 
        E => MSS_ADLIB_INST_MGPIO0B_OE, Y => GPIO_GPIO_0_BI_PAD_Y);
    
    FIC_2_APB_M_PCLK_inferred_clock_RNIPG5_0 : CFG1
      generic map(INIT => "01")

      port map(A => \CORECONFIGP_0_APB_S_PCLK\, Y => 
        CORECONFIGP_0_APB_S_PCLK_i);
    
    MDDR_ADDR_13_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[13]\, PAD => MDDR_ADDR(13));
    
    I2C_1_SDA_PAD : BIBUF
      port map(PAD => I2C_1_SDA, D => 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT, E => 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE, Y => 
        I2C_1_SDA_PAD_Y);
    
    I2C_1_SCL_PAD : BIBUF
      port map(PAD => I2C_1_SCL, D => 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT, E => 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE, Y => 
        I2C_1_SCL_PAD_Y);
    
    MDDR_ADDR_5_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[5]\, PAD => MDDR_ADDR(5));
    
    MDDR_DM_RDQS_1_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DM_RDQS(1), D => 
        \DRAM_DM_RDQS_OUT_net_0[1]\, E => \DM_OE_net_0[1]\, Y => 
        MDDR_DM_RDQS_1_PAD_Y);
    
    GPIO_GPIO_12_BI_PAD : BIBUF
      port map(PAD => GPIO_12_BI, D => 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OE, Y => 
        GPIO_GPIO_12_BI_PAD_Y);
    
    SPI_0_DO_PAD : TRIBUFF
      port map(D => MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        E => MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, PAD => 
        SPI_0_DO);
    
    MDDR_DQS_0_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQS(0), D => \DRAM_DQS_OUT_net_0[0]\, 
        E => \DRAM_DQS_OE_net_0[0]\, Y => MDDR_DQS_0_PAD_Y);
    
    MDDR_DQS_1_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQS(1), D => \DRAM_DQS_OUT_net_0[1]\, 
        E => \DRAM_DQS_OE_net_0[1]\, Y => MDDR_DQS_1_PAD_Y);
    
    MDDR_DQ_15_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(15), D => \DRAM_DQ_OUT_net_0[15]\, 
        E => \DRAM_DQ_OE_net_0[15]\, Y => MDDR_DQ_15_PAD_Y);
    
    MDDR_DM_RDQS_0_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DM_RDQS(0), D => 
        \DRAM_DM_RDQS_OUT_net_0[0]\, E => \DM_OE_net_0[0]\, Y => 
        MDDR_DM_RDQS_0_PAD_Y);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    SPI_0_DI_PAD : INBUF
      port map(PAD => SPI_0_DI, Y => SPI_0_DI_PAD_Y);
    
    MDDR_DQ_8_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(8), D => \DRAM_DQ_OUT_net_0[8]\, E
         => \DRAM_DQ_OE_net_0[8]\, Y => MDDR_DQ_8_PAD_Y);
    
    GPIO_GPIO_14_BI_PAD : BIBUF
      port map(PAD => GPIO_14_BI, D => 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OE, Y => 
        GPIO_GPIO_14_BI_PAD_Y);
    
    GPIO_GPIO_4_BI_PAD : BIBUF
      port map(PAD => GPIO_4_BI, D => 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT, E => 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE, Y => 
        GPIO_GPIO_4_BI_PAD_Y);
    
    MDDR_ADDR_9_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[9]\, PAD => MDDR_ADDR(9));
    
    MDDR_BA_2_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_BA_net_0[2]\, PAD => MDDR_BA(2));
    
    MDDR_ADDR_14_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[14]\, PAD => MDDR_ADDR(14));
    
    MSS_ADLIB_INST : MSS_060

              generic map(INIT => "00" & x"000000000000030000000000000003610008090A4290800908000000090A42000000000C03000000009000000000200012036190A4200001004000000000000000000000000000000000000F000000000000000000000000000000007FFFFFFFB000001007C35C804248006090801041A3FFFFE400000000000846809D001F0F41C00000002DA18010842108421000001FE34001FF8000000400000000020CD1007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
         ACT_UBITS => x"FFFFFFFFFFFFFF",
         MEMORYFILE => "ENVM_init.mem", RTC_MAIN_XTL_FREQ => 0.0,
         DDR_CLK_FREQ => 142.0)

      port map(CAN_RXBUS_MGPIO3A_H2F_A => OPEN, 
        CAN_RXBUS_MGPIO3A_H2F_B => OPEN, CAN_TX_EBL_MGPIO4A_H2F_A
         => OPEN, CAN_TX_EBL_MGPIO4A_H2F_B => OPEN, 
        CAN_TXBUS_MGPIO2A_H2F_A => OPEN, CAN_TXBUS_MGPIO2A_H2F_B
         => OPEN, CLK_CONFIG_APB => FIC_2_APB_M_PCLK, COMMS_INT
         => OPEN, CONFIG_PRESET_N => CONFIG_PRESET_N, 
        EDAC_ERROR(7) => nc228, EDAC_ERROR(6) => nc203, 
        EDAC_ERROR(5) => nc216, EDAC_ERROR(4) => nc194, 
        EDAC_ERROR(3) => nc151, EDAC_ERROR(2) => nc23, 
        EDAC_ERROR(1) => nc175, EDAC_ERROR(0) => nc58, 
        F_FM0_RDATA(31) => nc116, F_FM0_RDATA(30) => nc74, 
        F_FM0_RDATA(29) => nc133, F_FM0_RDATA(28) => nc238, 
        F_FM0_RDATA(27) => nc167, F_FM0_RDATA(26) => nc84, 
        F_FM0_RDATA(25) => nc39, F_FM0_RDATA(24) => nc72, 
        F_FM0_RDATA(23) => nc212, F_FM0_RDATA(22) => nc205, 
        F_FM0_RDATA(21) => nc82, F_FM0_RDATA(20) => nc145, 
        F_FM0_RDATA(19) => nc181, F_FM0_RDATA(18) => nc160, 
        F_FM0_RDATA(17) => nc57, F_FM0_RDATA(16) => nc156, 
        F_FM0_RDATA(15) => nc125, F_FM0_RDATA(14) => nc211, 
        F_FM0_RDATA(13) => nc73, F_FM0_RDATA(12) => nc107, 
        F_FM0_RDATA(11) => nc66, F_FM0_RDATA(10) => nc83, 
        F_FM0_RDATA(9) => nc9, F_FM0_RDATA(8) => nc171, 
        F_FM0_RDATA(7) => nc54, F_FM0_RDATA(6) => nc135, 
        F_FM0_RDATA(5) => nc41, F_FM0_RDATA(4) => nc100, 
        F_FM0_RDATA(3) => nc52, F_FM0_RDATA(2) => nc186, 
        F_FM0_RDATA(1) => nc29, F_FM0_RDATA(0) => nc118, 
        F_FM0_READYOUT => OPEN, F_FM0_RESP => OPEN, 
        F_HM0_ADDR(31) => nc60, F_HM0_ADDR(30) => nc141, 
        F_HM0_ADDR(29) => nc193, F_HM0_ADDR(28) => nc214, 
        F_HM0_ADDR(27) => nc240, F_HM0_ADDR(26) => nc45, 
        F_HM0_ADDR(25) => nc53, F_HM0_ADDR(24) => nc121, 
        F_HM0_ADDR(23) => nc176, F_HM0_ADDR(22) => nc220, 
        F_HM0_ADDR(21) => nc158, F_HM0_ADDR(20) => nc209, 
        F_HM0_ADDR(19) => nc246, F_HM0_ADDR(18) => nc162, 
        F_HM0_ADDR(17) => nc11, F_HM0_ADDR(16) => nc131, 
        F_HM0_ADDR(15) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15), 
        F_HM0_ADDR(14) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14), 
        F_HM0_ADDR(13) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13), 
        F_HM0_ADDR(12) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12), 
        F_HM0_ADDR(11) => nc96, F_HM0_ADDR(10) => nc79, 
        F_HM0_ADDR(9) => nc226, F_HM0_ADDR(8) => nc146, 
        F_HM0_ADDR(7) => CoreAPB3_0_APBmslave0_PADDR(7), 
        F_HM0_ADDR(6) => CoreAPB3_0_APBmslave0_PADDR(6), 
        F_HM0_ADDR(5) => CoreAPB3_0_APBmslave0_PADDR(5), 
        F_HM0_ADDR(4) => CoreAPB3_0_APBmslave0_PADDR(4), 
        F_HM0_ADDR(3) => CoreAPB3_0_APBmslave0_PADDR(3), 
        F_HM0_ADDR(2) => CoreAPB3_0_APBmslave0_PADDR(2), 
        F_HM0_ADDR(1) => CoreAPB3_0_APBmslave0_PADDR(1), 
        F_HM0_ADDR(0) => CoreAPB3_0_APBmslave0_PADDR(0), 
        F_HM0_ENABLE => CoreAPB3_0_APBmslave0_PENABLE, F_HM0_SEL
         => m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx, F_HM0_SIZE(1)
         => nc230, F_HM0_SIZE(0) => nc89, F_HM0_TRANS1 => OPEN, 
        F_HM0_WDATA(31) => nc119, F_HM0_WDATA(30) => nc48, 
        F_HM0_WDATA(29) => nc213, F_HM0_WDATA(28) => nc126, 
        F_HM0_WDATA(27) => nc195, F_HM0_WDATA(26) => nc188, 
        F_HM0_WDATA(25) => nc242, F_HM0_WDATA(24) => nc15, 
        F_HM0_WDATA(23) => nc236, F_HM0_WDATA(22) => nc102, 
        F_HM0_WDATA(21) => nc3, F_HM0_WDATA(20) => nc207, 
        F_HM0_WDATA(19) => nc47, F_HM0_WDATA(18) => nc90, 
        F_HM0_WDATA(17) => nc222, F_HM0_WDATA(16) => nc159, 
        F_HM0_WDATA(15) => nc136, F_HM0_WDATA(14) => nc241, 
        F_HM0_WDATA(13) => nc178, F_HM0_WDATA(12) => nc215, 
        F_HM0_WDATA(11) => nc59, F_HM0_WDATA(10) => nc221, 
        F_HM0_WDATA(9) => nc232, F_HM0_WDATA(8) => nc18, 
        F_HM0_WDATA(7) => CoreAPB3_0_APBmslave0_PWDATA(7), 
        F_HM0_WDATA(6) => CoreAPB3_0_APBmslave0_PWDATA(6), 
        F_HM0_WDATA(5) => CoreAPB3_0_APBmslave0_PWDATA(5), 
        F_HM0_WDATA(4) => CoreAPB3_0_APBmslave0_PWDATA(4), 
        F_HM0_WDATA(3) => CoreAPB3_0_APBmslave0_PWDATA(3), 
        F_HM0_WDATA(2) => CoreAPB3_0_APBmslave0_PWDATA(2), 
        F_HM0_WDATA(1) => CoreAPB3_0_APBmslave0_PWDATA(1), 
        F_HM0_WDATA(0) => CoreAPB3_0_APBmslave0_PWDATA(0), 
        F_HM0_WRITE => CoreAPB3_0_APBmslave0_PWRITE, FAB_CHRGVBUS
         => OPEN, FAB_DISCHRGVBUS => OPEN, FAB_DMPULLDOWN => OPEN, 
        FAB_DPPULLDOWN => OPEN, FAB_DRVVBUS => OPEN, FAB_IDPULLUP
         => OPEN, FAB_OPMODE(1) => nc44, FAB_OPMODE(0) => nc117, 
        FAB_SUSPENDM => OPEN, FAB_TERMSEL => OPEN, FAB_TXVALID
         => OPEN, FAB_VCONTROL(3) => nc189, FAB_VCONTROL(2) => 
        nc164, FAB_VCONTROL(1) => nc148, FAB_VCONTROL(0) => nc42, 
        FAB_VCONTROLLOADM => OPEN, FAB_XCVRSEL(1) => nc231, 
        FAB_XCVRSEL(0) => nc191, FAB_XDATAOUT(7) => nc17, 
        FAB_XDATAOUT(6) => nc2, FAB_XDATAOUT(5) => nc110, 
        FAB_XDATAOUT(4) => nc128, FAB_XDATAOUT(3) => nc244, 
        FAB_XDATAOUT(2) => nc43, FAB_XDATAOUT(1) => nc179, 
        FAB_XDATAOUT(0) => nc157, FACC_GLMUX_SEL => OPEN, 
        FIC32_0_MASTER(1) => nc36, FIC32_0_MASTER(0) => nc224, 
        FIC32_1_MASTER(1) => nc61, FIC32_1_MASTER(0) => nc104, 
        FPGA_RESET_N => m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        GTX_CLK => OPEN, H2F_INTERRUPT(15) => nc138, 
        H2F_INTERRUPT(14) => nc14, H2F_INTERRUPT(13) => nc150, 
        H2F_INTERRUPT(12) => nc196, H2F_INTERRUPT(11) => nc234, 
        H2F_INTERRUPT(10) => nc149, H2F_INTERRUPT(9) => nc12, 
        H2F_INTERRUPT(8) => nc219, H2F_INTERRUPT(7) => nc30, 
        H2F_INTERRUPT(6) => nc243, H2F_INTERRUPT(5) => nc187, 
        H2F_INTERRUPT(4) => nc65, H2F_INTERRUPT(3) => nc7, 
        H2F_INTERRUPT(2) => nc129, H2F_INTERRUPT(1) => nc8, 
        H2F_INTERRUPT(0) => nc223, H2F_NMI => OPEN, H2FCALIB => 
        OPEN, I2C0_SCL_MGPIO31B_H2F_A => OPEN, 
        I2C0_SCL_MGPIO31B_H2F_B => OPEN, I2C0_SDA_MGPIO30B_H2F_A
         => OPEN, I2C0_SDA_MGPIO30B_H2F_B => OPEN, 
        I2C1_SCL_MGPIO1A_H2F_A => 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE, I2C1_SCL_MGPIO1A_H2F_B
         => GPIO_1_M2F, I2C1_SDA_MGPIO0A_H2F_A => OPEN, 
        I2C1_SDA_MGPIO0A_H2F_B => OPEN, MDCF => MAC_MII_MDC_c, 
        MDOENF => m2s010_som_sb_MSS_0_MAC_MII_MDO_EN, MDOF => 
        m2s010_som_sb_MSS_0_MAC_MII_MDO, 
        MMUART0_CTS_MGPIO19B_H2F_A => OPEN, 
        MMUART0_CTS_MGPIO19B_H2F_B => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_A => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_B => GPIO_22_M2F_c, 
        MMUART0_DSR_MGPIO20B_H2F_A => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_B => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_A => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_B => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_A => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_B => GPIO_21_M2F_c, 
        MMUART0_RTS_MGPIO17B_H2F_A => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_B => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_A => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_B => 
        m2s010_som_sb_0_GPIO_28_SW_RESET, 
        MMUART0_SCK_MGPIO29B_H2F_A => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_B => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_A => MMUART_0_TXD_M2F_c, 
        MMUART0_TXD_MGPIO27B_H2F_B => OPEN, 
        MMUART1_DTR_MGPIO12B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_B => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_A => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_B => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_A => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_B => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_A => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_B => GPIO_24_M2F_c, MPLL_LOCK
         => OPEN, PER2_FABRIC_PADDR(15) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(15), 
        PER2_FABRIC_PADDR(14) => nc13, PER2_FABRIC_PADDR(13) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(13), 
        PER2_FABRIC_PADDR(12) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(12), 
        PER2_FABRIC_PADDR(11) => nc180, PER2_FABRIC_PADDR(10) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(10), 
        PER2_FABRIC_PADDR(9) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(9), 
        PER2_FABRIC_PADDR(8) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(8), 
        PER2_FABRIC_PADDR(7) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(7), 
        PER2_FABRIC_PADDR(6) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(6), 
        PER2_FABRIC_PADDR(5) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(5), 
        PER2_FABRIC_PADDR(4) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), 
        PER2_FABRIC_PADDR(3) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), 
        PER2_FABRIC_PADDR(2) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), 
        PER2_FABRIC_PENABLE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, 
        PER2_FABRIC_PSEL => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx, 
        PER2_FABRIC_PWDATA(31) => nc26, PER2_FABRIC_PWDATA(30)
         => nc177, PER2_FABRIC_PWDATA(29) => nc139, 
        PER2_FABRIC_PWDATA(28) => nc245, PER2_FABRIC_PWDATA(27)
         => nc233, PER2_FABRIC_PWDATA(26) => nc163, 
        PER2_FABRIC_PWDATA(25) => nc112, PER2_FABRIC_PWDATA(24)
         => nc68, PER2_FABRIC_PWDATA(23) => nc49, 
        PER2_FABRIC_PWDATA(22) => nc217, PER2_FABRIC_PWDATA(21)
         => nc170, PER2_FABRIC_PWDATA(20) => nc91, 
        PER2_FABRIC_PWDATA(19) => nc225, PER2_FABRIC_PWDATA(18)
         => nc5, PER2_FABRIC_PWDATA(17) => nc20, 
        PER2_FABRIC_PWDATA(16) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(16), 
        PER2_FABRIC_PWDATA(15) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(15), 
        PER2_FABRIC_PWDATA(14) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(14), 
        PER2_FABRIC_PWDATA(13) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(13), 
        PER2_FABRIC_PWDATA(12) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(12), 
        PER2_FABRIC_PWDATA(11) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(11), 
        PER2_FABRIC_PWDATA(10) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(10), 
        PER2_FABRIC_PWDATA(9) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(9), 
        PER2_FABRIC_PWDATA(8) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(8), 
        PER2_FABRIC_PWDATA(7) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(7), 
        PER2_FABRIC_PWDATA(6) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(6), 
        PER2_FABRIC_PWDATA(5) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(5), 
        PER2_FABRIC_PWDATA(4) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(4), 
        PER2_FABRIC_PWDATA(3) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(3), 
        PER2_FABRIC_PWDATA(2) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(2), 
        PER2_FABRIC_PWDATA(1) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1), 
        PER2_FABRIC_PWDATA(0) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0), 
        PER2_FABRIC_PWRITE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, 
        RTC_MATCH => OPEN, SLEEPDEEP => OPEN, SLEEPHOLDACK => 
        OPEN, SLEEPING => OPEN, SMBALERT_NO0 => OPEN, 
        SMBALERT_NO1 => OPEN, SMBSUS_NO0 => OPEN, SMBSUS_NO1 => 
        OPEN, SPI0_CLK_OUT => OPEN, SPI0_SDI_MGPIO5A_H2F_A => 
        OPEN, SPI0_SDI_MGPIO5A_H2F_B => GPIO_5_M2F_c, 
        SPI0_SDO_MGPIO6A_H2F_A => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F_OE, SPI0_SDO_MGPIO6A_H2F_B
         => m2s010_som_sb_MSS_0_GPIO_6_M2F, 
        SPI0_SS0_MGPIO7A_H2F_A => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE, SPI0_SS0_MGPIO7A_H2F_B
         => m2s010_som_sb_MSS_0_GPIO_7_M2F, 
        SPI0_SS1_MGPIO8A_H2F_A => OPEN, SPI0_SS1_MGPIO8A_H2F_B
         => GPIO_8_M2F_c, SPI0_SS2_MGPIO9A_H2F_A => OPEN, 
        SPI0_SS2_MGPIO9A_H2F_B => OPEN, SPI0_SS3_MGPIO10A_H2F_A
         => OPEN, SPI0_SS3_MGPIO10A_H2F_B => OPEN, 
        SPI0_SS4_MGPIO19A_H2F_A => OPEN, SPI0_SS5_MGPIO20A_H2F_A
         => OPEN, SPI0_SS6_MGPIO21A_H2F_A => OPEN, 
        SPI0_SS7_MGPIO22A_H2F_A => OPEN, SPI1_CLK_OUT => 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F, 
        SPI1_SDI_MGPIO11A_H2F_A => OPEN, SPI1_SDI_MGPIO11A_H2F_B
         => GPIO_11_M2F_c, SPI1_SDO_MGPIO12A_H2F_A => 
        SPI_1_DO_CAM_c, SPI1_SDO_MGPIO12A_H2F_B => OPEN, 
        SPI1_SS0_MGPIO13A_H2F_A => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F, 
        SPI1_SS0_MGPIO13A_H2F_B => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        SPI1_SS1_MGPIO14A_H2F_A => OPEN, SPI1_SS1_MGPIO14A_H2F_B
         => OPEN, SPI1_SS2_MGPIO15A_H2F_A => OPEN, 
        SPI1_SS2_MGPIO15A_H2F_B => OPEN, SPI1_SS3_MGPIO16A_H2F_A
         => OPEN, SPI1_SS3_MGPIO16A_H2F_B => OPEN, 
        SPI1_SS4_MGPIO17A_H2F_A => OPEN, SPI1_SS5_MGPIO18A_H2F_A
         => OPEN, SPI1_SS6_MGPIO23A_H2F_A => OPEN, 
        SPI1_SS7_MGPIO24A_H2F_A => OPEN, TCGF(9) => nc198, 
        TCGF(8) => nc147, TCGF(7) => nc67, TCGF(6) => nc152, 
        TCGF(5) => nc127, TCGF(4) => nc103, TCGF(3) => nc235, 
        TCGF(2) => nc76, TCGF(1) => nc208, TCGF(0) => nc140, 
        TRACECLK => OPEN, TRACEDATA(3) => nc86, TRACEDATA(2) => 
        nc95, TRACEDATA(1) => nc120, TRACEDATA(0) => nc165, 
        TX_CLK => OPEN, TX_ENF => MAC_MII_TX_EN_c, TX_ERRF => 
        OPEN, TXCTL_EN_RIF => OPEN, TXD_RIF(3) => nc137, 
        TXD_RIF(2) => nc64, TXD_RIF(1) => nc19, TXD_RIF(0) => 
        nc70, TXDF(7) => nc182, TXDF(6) => nc62, TXDF(5) => nc199, 
        TXDF(4) => nc80, TXDF(3) => MAC_MII_TXD_c(3), TXDF(2) => 
        MAC_MII_TXD_c(2), TXDF(1) => MAC_MII_TXD_c(1), TXDF(0)
         => MAC_MII_TXD_c(0), TXEV => OPEN, WDOGTIMEOUT => OPEN, 
        F_ARREADY_HREADYOUT1 => OPEN, F_AWREADY_HREADYOUT0 => 
        OPEN, F_BID(3) => nc130, F_BID(2) => nc98, F_BID(1) => 
        nc114, F_BID(0) => nc56, F_BRESP_HRESP0(1) => nc105, 
        F_BRESP_HRESP0(0) => nc63, F_BVALID => OPEN, 
        F_RDATA_HRDATA01(63) => nc172, F_RDATA_HRDATA01(62) => 
        nc229, F_RDATA_HRDATA01(61) => nc97, F_RDATA_HRDATA01(60)
         => nc161, F_RDATA_HRDATA01(59) => nc31, 
        F_RDATA_HRDATA01(58) => nc154, F_RDATA_HRDATA01(57) => 
        nc50, F_RDATA_HRDATA01(56) => nc239, F_RDATA_HRDATA01(55)
         => nc142, F_RDATA_HRDATA01(54) => nc94, 
        F_RDATA_HRDATA01(53) => nc197, F_RDATA_HRDATA01(52) => 
        nc122, F_RDATA_HRDATA01(51) => nc35, F_RDATA_HRDATA01(50)
         => nc4, F_RDATA_HRDATA01(49) => nc227, 
        F_RDATA_HRDATA01(48) => nc92, F_RDATA_HRDATA01(47) => 
        nc101, F_RDATA_HRDATA01(46) => nc184, 
        F_RDATA_HRDATA01(45) => nc200, F_RDATA_HRDATA01(44) => 
        nc190, F_RDATA_HRDATA01(43) => nc166, 
        F_RDATA_HRDATA01(42) => nc132, F_RDATA_HRDATA01(41) => 
        nc21, F_RDATA_HRDATA01(40) => nc237, F_RDATA_HRDATA01(39)
         => nc93, F_RDATA_HRDATA01(38) => nc69, 
        F_RDATA_HRDATA01(37) => nc206, F_RDATA_HRDATA01(36) => 
        nc174, F_RDATA_HRDATA01(35) => nc38, F_RDATA_HRDATA01(34)
         => nc113, F_RDATA_HRDATA01(33) => nc218, 
        F_RDATA_HRDATA01(32) => nc106, F_RDATA_HRDATA01(31) => 
        nc25, F_RDATA_HRDATA01(30) => nc1, F_RDATA_HRDATA01(29)
         => nc37, F_RDATA_HRDATA01(28) => nc202, 
        F_RDATA_HRDATA01(27) => nc144, F_RDATA_HRDATA01(26) => 
        nc153, F_RDATA_HRDATA01(25) => nc46, F_RDATA_HRDATA01(24)
         => nc71, F_RDATA_HRDATA01(23) => nc124, 
        F_RDATA_HRDATA01(22) => nc81, F_RDATA_HRDATA01(21) => 
        nc201, F_RDATA_HRDATA01(20) => nc168, 
        F_RDATA_HRDATA01(19) => nc34, F_RDATA_HRDATA01(18) => 
        nc28, F_RDATA_HRDATA01(17) => nc115, F_RDATA_HRDATA01(16)
         => nc192, F_RDATA_HRDATA01(15) => nc134, 
        F_RDATA_HRDATA01(14) => nc32, F_RDATA_HRDATA01(13) => 
        nc40, F_RDATA_HRDATA01(12) => nc99, F_RDATA_HRDATA01(11)
         => nc75, F_RDATA_HRDATA01(10) => nc183, 
        F_RDATA_HRDATA01(9) => nc85, F_RDATA_HRDATA01(8) => nc27, 
        F_RDATA_HRDATA01(7) => nc108, F_RDATA_HRDATA01(6) => nc16, 
        F_RDATA_HRDATA01(5) => nc155, F_RDATA_HRDATA01(4) => nc51, 
        F_RDATA_HRDATA01(3) => nc33, F_RDATA_HRDATA01(2) => nc204, 
        F_RDATA_HRDATA01(1) => nc173, F_RDATA_HRDATA01(0) => 
        nc169, F_RID(3) => nc78, F_RID(2) => nc24, F_RID(1) => 
        nc88, F_RID(0) => nc111, F_RLAST => OPEN, 
        F_RRESP_HRESP1(1) => nc55, F_RRESP_HRESP1(0) => nc10, 
        F_RVALID => OPEN, F_WREADY => OPEN, 
        MDDR_FABRIC_PRDATA(15) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(15), 
        MDDR_FABRIC_PRDATA(14) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(14), 
        MDDR_FABRIC_PRDATA(13) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(13), 
        MDDR_FABRIC_PRDATA(12) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(12), 
        MDDR_FABRIC_PRDATA(11) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(11), 
        MDDR_FABRIC_PRDATA(10) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(10), 
        MDDR_FABRIC_PRDATA(9) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(9), 
        MDDR_FABRIC_PRDATA(8) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(8), 
        MDDR_FABRIC_PRDATA(7) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(7), 
        MDDR_FABRIC_PRDATA(6) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(6), 
        MDDR_FABRIC_PRDATA(5) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(5), 
        MDDR_FABRIC_PRDATA(4) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(4), 
        MDDR_FABRIC_PRDATA(3) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(3), 
        MDDR_FABRIC_PRDATA(2) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(2), 
        MDDR_FABRIC_PRDATA(1) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(1), 
        MDDR_FABRIC_PRDATA(0) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(0), 
        MDDR_FABRIC_PREADY => CORECONFIGP_0_MDDR_APBmslave_PREADY, 
        MDDR_FABRIC_PSLVERR => 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR, CAN_RXBUS_F2H_SCP
         => VCC_net_1, CAN_TX_EBL_F2H_SCP => VCC_net_1, 
        CAN_TXBUS_F2H_SCP => VCC_net_1, COLF => MAC_MII_COL_c, 
        CRSF => MAC_MII_CRS_c, F2_DMAREADY(1) => VCC_net_1, 
        F2_DMAREADY(0) => VCC_net_1, F2H_INTERRUPT(15) => 
        GND_net_1, F2H_INTERRUPT(14) => GND_net_1, 
        F2H_INTERRUPT(13) => GND_net_1, F2H_INTERRUPT(12) => 
        GND_net_1, F2H_INTERRUPT(11) => GND_net_1, 
        F2H_INTERRUPT(10) => GND_net_1, F2H_INTERRUPT(9) => 
        GND_net_1, F2H_INTERRUPT(8) => GND_net_1, 
        F2H_INTERRUPT(7) => GND_net_1, F2H_INTERRUPT(6) => 
        GND_net_1, F2H_INTERRUPT(5) => GND_net_1, 
        F2H_INTERRUPT(4) => GND_net_1, F2H_INTERRUPT(3) => 
        GND_net_1, F2H_INTERRUPT(2) => GND_net_1, 
        F2H_INTERRUPT(1) => GND_net_1, F2H_INTERRUPT(0) => 
        CommsFPGA_top_0_INT, F2HCALIB => VCC_net_1, F_DMAREADY(1)
         => VCC_net_1, F_DMAREADY(0) => VCC_net_1, F_FM0_ADDR(31)
         => GND_net_1, F_FM0_ADDR(30) => GND_net_1, 
        F_FM0_ADDR(29) => GND_net_1, F_FM0_ADDR(28) => GND_net_1, 
        F_FM0_ADDR(27) => GND_net_1, F_FM0_ADDR(26) => GND_net_1, 
        F_FM0_ADDR(25) => GND_net_1, F_FM0_ADDR(24) => GND_net_1, 
        F_FM0_ADDR(23) => GND_net_1, F_FM0_ADDR(22) => GND_net_1, 
        F_FM0_ADDR(21) => GND_net_1, F_FM0_ADDR(20) => GND_net_1, 
        F_FM0_ADDR(19) => GND_net_1, F_FM0_ADDR(18) => GND_net_1, 
        F_FM0_ADDR(17) => GND_net_1, F_FM0_ADDR(16) => GND_net_1, 
        F_FM0_ADDR(15) => GND_net_1, F_FM0_ADDR(14) => GND_net_1, 
        F_FM0_ADDR(13) => GND_net_1, F_FM0_ADDR(12) => GND_net_1, 
        F_FM0_ADDR(11) => GND_net_1, F_FM0_ADDR(10) => GND_net_1, 
        F_FM0_ADDR(9) => GND_net_1, F_FM0_ADDR(8) => GND_net_1, 
        F_FM0_ADDR(7) => GND_net_1, F_FM0_ADDR(6) => GND_net_1, 
        F_FM0_ADDR(5) => GND_net_1, F_FM0_ADDR(4) => GND_net_1, 
        F_FM0_ADDR(3) => GND_net_1, F_FM0_ADDR(2) => GND_net_1, 
        F_FM0_ADDR(1) => GND_net_1, F_FM0_ADDR(0) => GND_net_1, 
        F_FM0_ENABLE => GND_net_1, F_FM0_MASTLOCK => GND_net_1, 
        F_FM0_READY => VCC_net_1, F_FM0_SEL => GND_net_1, 
        F_FM0_SIZE(1) => GND_net_1, F_FM0_SIZE(0) => GND_net_1, 
        F_FM0_TRANS1 => GND_net_1, F_FM0_WDATA(31) => GND_net_1, 
        F_FM0_WDATA(30) => GND_net_1, F_FM0_WDATA(29) => 
        GND_net_1, F_FM0_WDATA(28) => GND_net_1, F_FM0_WDATA(27)
         => GND_net_1, F_FM0_WDATA(26) => GND_net_1, 
        F_FM0_WDATA(25) => GND_net_1, F_FM0_WDATA(24) => 
        GND_net_1, F_FM0_WDATA(23) => GND_net_1, F_FM0_WDATA(22)
         => GND_net_1, F_FM0_WDATA(21) => GND_net_1, 
        F_FM0_WDATA(20) => GND_net_1, F_FM0_WDATA(19) => 
        GND_net_1, F_FM0_WDATA(18) => GND_net_1, F_FM0_WDATA(17)
         => GND_net_1, F_FM0_WDATA(16) => GND_net_1, 
        F_FM0_WDATA(15) => GND_net_1, F_FM0_WDATA(14) => 
        GND_net_1, F_FM0_WDATA(13) => GND_net_1, F_FM0_WDATA(12)
         => GND_net_1, F_FM0_WDATA(11) => GND_net_1, 
        F_FM0_WDATA(10) => GND_net_1, F_FM0_WDATA(9) => GND_net_1, 
        F_FM0_WDATA(8) => GND_net_1, F_FM0_WDATA(7) => GND_net_1, 
        F_FM0_WDATA(6) => GND_net_1, F_FM0_WDATA(5) => GND_net_1, 
        F_FM0_WDATA(4) => GND_net_1, F_FM0_WDATA(3) => GND_net_1, 
        F_FM0_WDATA(2) => GND_net_1, F_FM0_WDATA(1) => GND_net_1, 
        F_FM0_WDATA(0) => GND_net_1, F_FM0_WRITE => GND_net_1, 
        F_HM0_RDATA(31) => GND_net_1, F_HM0_RDATA(30) => 
        GND_net_1, F_HM0_RDATA(29) => GND_net_1, F_HM0_RDATA(28)
         => GND_net_1, F_HM0_RDATA(27) => GND_net_1, 
        F_HM0_RDATA(26) => GND_net_1, F_HM0_RDATA(25) => 
        GND_net_1, F_HM0_RDATA(24) => GND_net_1, F_HM0_RDATA(23)
         => GND_net_1, F_HM0_RDATA(22) => GND_net_1, 
        F_HM0_RDATA(21) => GND_net_1, F_HM0_RDATA(20) => 
        GND_net_1, F_HM0_RDATA(19) => GND_net_1, F_HM0_RDATA(18)
         => GND_net_1, F_HM0_RDATA(17) => GND_net_1, 
        F_HM0_RDATA(16) => GND_net_1, F_HM0_RDATA(15) => 
        GND_net_1, F_HM0_RDATA(14) => GND_net_1, F_HM0_RDATA(13)
         => GND_net_1, F_HM0_RDATA(12) => GND_net_1, 
        F_HM0_RDATA(11) => GND_net_1, F_HM0_RDATA(10) => 
        GND_net_1, F_HM0_RDATA(9) => GND_net_1, F_HM0_RDATA(8)
         => GND_net_1, F_HM0_RDATA(7) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(7), F_HM0_RDATA(6) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(6), F_HM0_RDATA(5) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(5), F_HM0_RDATA(4) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(4), F_HM0_RDATA(3) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(3), F_HM0_RDATA(2) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(2), F_HM0_RDATA(1) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(1), F_HM0_RDATA(0) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(0), F_HM0_READY => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, F_HM0_RESP => 
        GND_net_1, FAB_AVALID => VCC_net_1, FAB_HOSTDISCON => 
        VCC_net_1, FAB_IDDIG => VCC_net_1, FAB_LINESTATE(1) => 
        VCC_net_1, FAB_LINESTATE(0) => VCC_net_1, FAB_M3_RESET_N
         => VCC_net_1, FAB_PLL_LOCK => FAB_CCC_LOCK, FAB_RXACTIVE
         => VCC_net_1, FAB_RXERROR => VCC_net_1, FAB_RXVALID => 
        VCC_net_1, FAB_RXVALIDH => GND_net_1, FAB_SESSEND => 
        VCC_net_1, FAB_TXREADY => VCC_net_1, FAB_VBUSVALID => 
        VCC_net_1, FAB_VSTATUS(7) => VCC_net_1, FAB_VSTATUS(6)
         => VCC_net_1, FAB_VSTATUS(5) => VCC_net_1, 
        FAB_VSTATUS(4) => VCC_net_1, FAB_VSTATUS(3) => VCC_net_1, 
        FAB_VSTATUS(2) => VCC_net_1, FAB_VSTATUS(1) => VCC_net_1, 
        FAB_VSTATUS(0) => VCC_net_1, FAB_XDATAIN(7) => VCC_net_1, 
        FAB_XDATAIN(6) => VCC_net_1, FAB_XDATAIN(5) => VCC_net_1, 
        FAB_XDATAIN(4) => VCC_net_1, FAB_XDATAIN(3) => VCC_net_1, 
        FAB_XDATAIN(2) => VCC_net_1, FAB_XDATAIN(1) => VCC_net_1, 
        FAB_XDATAIN(0) => VCC_net_1, GTX_CLKPF => VCC_net_1, 
        I2C0_BCLK => VCC_net_1, I2C0_SCL_F2H_SCP => VCC_net_1, 
        I2C0_SDA_F2H_SCP => VCC_net_1, I2C1_BCLK => VCC_net_1, 
        I2C1_SCL_F2H_SCP => VCC_net_1, I2C1_SDA_F2H_SCP => 
        VCC_net_1, MDIF => BIBUF_0_Y, MGPIO0A_F2H_GPIN => 
        VCC_net_1, MGPIO10A_F2H_GPIN => Y_net_0(3), 
        MGPIO11A_F2H_GPIN => VCC_net_1, MGPIO11B_F2H_GPIN => 
        VCC_net_1, MGPIO12A_F2H_GPIN => VCC_net_1, 
        MGPIO13A_F2H_GPIN => VCC_net_1, MGPIO14A_F2H_GPIN => 
        VCC_net_1, MGPIO15A_F2H_GPIN => VCC_net_1, 
        MGPIO16A_F2H_GPIN => VCC_net_1, MGPIO17B_F2H_GPIN => 
        VCC_net_1, MGPIO18B_F2H_GPIN => VCC_net_1, 
        MGPIO19B_F2H_GPIN => Y_net_0(1), MGPIO1A_F2H_GPIN => 
        GPIO_1_in_0, MGPIO20B_F2H_GPIN => VCC_net_1, 
        MGPIO21B_F2H_GPIN => VCC_net_1, MGPIO22B_F2H_GPIN => 
        VCC_net_1, MGPIO24B_F2H_GPIN => VCC_net_1, 
        MGPIO25B_F2H_GPIN => VCC_net_1, MGPIO26B_F2H_GPIN => 
        VCC_net_1, MGPIO27B_F2H_GPIN => DEBOUNCE_OUT_1_c, 
        MGPIO28B_F2H_GPIN => VCC_net_1, MGPIO29B_F2H_GPIN => 
        DEBOUNCE_OUT_2_c, MGPIO2A_F2H_GPIN => Y_net_0(2), 
        MGPIO30B_F2H_GPIN => DEBOUNCE_OUT_net_0_0, 
        MGPIO31B_F2H_GPIN => VCC_net_1, MGPIO3A_F2H_GPIN => 
        VCC_net_1, MGPIO4A_F2H_GPIN => VCC_net_1, 
        MGPIO5A_F2H_GPIN => VCC_net_1, MGPIO6A_F2H_GPIN => 
        GPIO_6_Y_0, MGPIO7A_F2H_GPIN => GPIO_7_Y_0, 
        MGPIO8A_F2H_GPIN => VCC_net_1, MGPIO9A_F2H_GPIN => 
        Y_net_0(0), MMUART0_CTS_F2H_SCP => VCC_net_1, 
        MMUART0_DCD_F2H_SCP => VCC_net_1, MMUART0_DSR_F2H_SCP => 
        VCC_net_1, MMUART0_DTR_F2H_SCP => VCC_net_1, 
        MMUART0_RI_F2H_SCP => VCC_net_1, MMUART0_RTS_F2H_SCP => 
        VCC_net_1, MMUART0_RXD_F2H_SCP => MMUART_0_RXD_F2M_c, 
        MMUART0_SCK_F2H_SCP => VCC_net_1, MMUART0_TXD_F2H_SCP => 
        VCC_net_1, MMUART1_CTS_F2H_SCP => VCC_net_1, 
        MMUART1_DCD_F2H_SCP => VCC_net_1, MMUART1_DSR_F2H_SCP => 
        VCC_net_1, MMUART1_RI_F2H_SCP => VCC_net_1, 
        MMUART1_RTS_F2H_SCP => VCC_net_1, MMUART1_RXD_F2H_SCP => 
        VCC_net_1, MMUART1_SCK_F2H_SCP => VCC_net_1, 
        MMUART1_TXD_F2H_SCP => VCC_net_1, PER2_FABRIC_PRDATA(31)
         => GND_net_1, PER2_FABRIC_PRDATA(30) => GND_net_1, 
        PER2_FABRIC_PRDATA(29) => GND_net_1, 
        PER2_FABRIC_PRDATA(28) => GND_net_1, 
        PER2_FABRIC_PRDATA(27) => GND_net_1, 
        PER2_FABRIC_PRDATA(26) => GND_net_1, 
        PER2_FABRIC_PRDATA(25) => GND_net_1, 
        PER2_FABRIC_PRDATA(24) => GND_net_1, 
        PER2_FABRIC_PRDATA(23) => GND_net_1, 
        PER2_FABRIC_PRDATA(22) => GND_net_1, 
        PER2_FABRIC_PRDATA(21) => GND_net_1, 
        PER2_FABRIC_PRDATA(20) => GND_net_1, 
        PER2_FABRIC_PRDATA(19) => GND_net_1, 
        PER2_FABRIC_PRDATA(18) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(17), 
        PER2_FABRIC_PRDATA(17) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(17), 
        PER2_FABRIC_PRDATA(16) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(16), 
        PER2_FABRIC_PRDATA(15) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(15), 
        PER2_FABRIC_PRDATA(14) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(14), 
        PER2_FABRIC_PRDATA(13) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(13), 
        PER2_FABRIC_PRDATA(12) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(12), 
        PER2_FABRIC_PRDATA(11) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(11), 
        PER2_FABRIC_PRDATA(10) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(10), 
        PER2_FABRIC_PRDATA(9) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(9), 
        PER2_FABRIC_PRDATA(8) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(8), 
        PER2_FABRIC_PRDATA(7) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(7), 
        PER2_FABRIC_PRDATA(6) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(6), 
        PER2_FABRIC_PRDATA(5) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(5), 
        PER2_FABRIC_PRDATA(4) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(4), 
        PER2_FABRIC_PRDATA(3) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(3), 
        PER2_FABRIC_PRDATA(2) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(2), 
        PER2_FABRIC_PRDATA(1) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(1), 
        PER2_FABRIC_PRDATA(0) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(0), 
        PER2_FABRIC_PREADY => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY, 
        PER2_FABRIC_PSLVERR => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR, RCGF(9)
         => VCC_net_1, RCGF(8) => VCC_net_1, RCGF(7) => VCC_net_1, 
        RCGF(6) => VCC_net_1, RCGF(5) => VCC_net_1, RCGF(4) => 
        VCC_net_1, RCGF(3) => VCC_net_1, RCGF(2) => VCC_net_1, 
        RCGF(1) => VCC_net_1, RCGF(0) => VCC_net_1, RX_CLKPF => 
        MAC_MII_RX_CLK_c, RX_DVF => MAC_MII_RX_DV_c, RX_ERRF => 
        MAC_MII_RX_ER_c, RX_EV => VCC_net_1, RXDF(7) => VCC_net_1, 
        RXDF(6) => VCC_net_1, RXDF(5) => VCC_net_1, RXDF(4) => 
        VCC_net_1, RXDF(3) => MAC_MII_RXD_c(3), RXDF(2) => 
        MAC_MII_RXD_c(2), RXDF(1) => MAC_MII_RXD_c(1), RXDF(0)
         => MAC_MII_RXD_c(0), SLEEPHOLDREQ => GND_net_1, 
        SMBALERT_NI0 => VCC_net_1, SMBALERT_NI1 => VCC_net_1, 
        SMBSUS_NI0 => VCC_net_1, SMBSUS_NI1 => VCC_net_1, 
        SPI0_CLK_IN => VCC_net_1, SPI0_SDI_F2H_SCP => VCC_net_1, 
        SPI0_SDO_F2H_SCP => VCC_net_1, SPI0_SS0_F2H_SCP => 
        VCC_net_1, SPI0_SS1_F2H_SCP => VCC_net_1, 
        SPI0_SS2_F2H_SCP => VCC_net_1, SPI0_SS3_F2H_SCP => 
        VCC_net_1, SPI1_CLK_IN => CAM_SPI_1_CLK_Y_0, 
        SPI1_SDI_F2H_SCP => SPI_1_DI, SPI1_SDO_F2H_SCP => 
        VCC_net_1, SPI1_SS0_F2H_SCP => SPI_1_SS0_MX_Y, 
        SPI1_SS1_F2H_SCP => VCC_net_1, SPI1_SS2_F2H_SCP => 
        VCC_net_1, SPI1_SS3_F2H_SCP => VCC_net_1, TX_CLKPF => 
        MAC_MII_TX_CLK_c, USER_MSS_GPIO_RESET_N => VCC_net_1, 
        USER_MSS_RESET_N => VCC_net_1, XCLK_FAB => VCC_net_1, 
        CLK_BASE => m2s010_som_sb_0_CCC_71MHz, CLK_MDDR_APB => 
        \CORECONFIGP_0_APB_S_PCLK\, F_ARADDR_HADDR1(31) => 
        VCC_net_1, F_ARADDR_HADDR1(30) => VCC_net_1, 
        F_ARADDR_HADDR1(29) => VCC_net_1, F_ARADDR_HADDR1(28) => 
        VCC_net_1, F_ARADDR_HADDR1(27) => VCC_net_1, 
        F_ARADDR_HADDR1(26) => VCC_net_1, F_ARADDR_HADDR1(25) => 
        VCC_net_1, F_ARADDR_HADDR1(24) => VCC_net_1, 
        F_ARADDR_HADDR1(23) => VCC_net_1, F_ARADDR_HADDR1(22) => 
        VCC_net_1, F_ARADDR_HADDR1(21) => VCC_net_1, 
        F_ARADDR_HADDR1(20) => VCC_net_1, F_ARADDR_HADDR1(19) => 
        VCC_net_1, F_ARADDR_HADDR1(18) => VCC_net_1, 
        F_ARADDR_HADDR1(17) => VCC_net_1, F_ARADDR_HADDR1(16) => 
        VCC_net_1, F_ARADDR_HADDR1(15) => VCC_net_1, 
        F_ARADDR_HADDR1(14) => VCC_net_1, F_ARADDR_HADDR1(13) => 
        VCC_net_1, F_ARADDR_HADDR1(12) => VCC_net_1, 
        F_ARADDR_HADDR1(11) => VCC_net_1, F_ARADDR_HADDR1(10) => 
        VCC_net_1, F_ARADDR_HADDR1(9) => VCC_net_1, 
        F_ARADDR_HADDR1(8) => VCC_net_1, F_ARADDR_HADDR1(7) => 
        VCC_net_1, F_ARADDR_HADDR1(6) => VCC_net_1, 
        F_ARADDR_HADDR1(5) => VCC_net_1, F_ARADDR_HADDR1(4) => 
        VCC_net_1, F_ARADDR_HADDR1(3) => VCC_net_1, 
        F_ARADDR_HADDR1(2) => VCC_net_1, F_ARADDR_HADDR1(1) => 
        VCC_net_1, F_ARADDR_HADDR1(0) => VCC_net_1, 
        F_ARBURST_HTRANS1(1) => GND_net_1, F_ARBURST_HTRANS1(0)
         => GND_net_1, F_ARID_HSEL1(3) => GND_net_1, 
        F_ARID_HSEL1(2) => GND_net_1, F_ARID_HSEL1(1) => 
        GND_net_1, F_ARID_HSEL1(0) => GND_net_1, 
        F_ARLEN_HBURST1(3) => GND_net_1, F_ARLEN_HBURST1(2) => 
        GND_net_1, F_ARLEN_HBURST1(1) => GND_net_1, 
        F_ARLEN_HBURST1(0) => GND_net_1, F_ARLOCK_HMASTLOCK1(1)
         => GND_net_1, F_ARLOCK_HMASTLOCK1(0) => GND_net_1, 
        F_ARSIZE_HSIZE1(1) => GND_net_1, F_ARSIZE_HSIZE1(0) => 
        GND_net_1, F_ARVALID_HWRITE1 => GND_net_1, 
        F_AWADDR_HADDR0(31) => VCC_net_1, F_AWADDR_HADDR0(30) => 
        VCC_net_1, F_AWADDR_HADDR0(29) => VCC_net_1, 
        F_AWADDR_HADDR0(28) => VCC_net_1, F_AWADDR_HADDR0(27) => 
        VCC_net_1, F_AWADDR_HADDR0(26) => VCC_net_1, 
        F_AWADDR_HADDR0(25) => VCC_net_1, F_AWADDR_HADDR0(24) => 
        VCC_net_1, F_AWADDR_HADDR0(23) => VCC_net_1, 
        F_AWADDR_HADDR0(22) => VCC_net_1, F_AWADDR_HADDR0(21) => 
        VCC_net_1, F_AWADDR_HADDR0(20) => VCC_net_1, 
        F_AWADDR_HADDR0(19) => VCC_net_1, F_AWADDR_HADDR0(18) => 
        VCC_net_1, F_AWADDR_HADDR0(17) => VCC_net_1, 
        F_AWADDR_HADDR0(16) => VCC_net_1, F_AWADDR_HADDR0(15) => 
        VCC_net_1, F_AWADDR_HADDR0(14) => VCC_net_1, 
        F_AWADDR_HADDR0(13) => VCC_net_1, F_AWADDR_HADDR0(12) => 
        VCC_net_1, F_AWADDR_HADDR0(11) => VCC_net_1, 
        F_AWADDR_HADDR0(10) => VCC_net_1, F_AWADDR_HADDR0(9) => 
        VCC_net_1, F_AWADDR_HADDR0(8) => VCC_net_1, 
        F_AWADDR_HADDR0(7) => VCC_net_1, F_AWADDR_HADDR0(6) => 
        VCC_net_1, F_AWADDR_HADDR0(5) => VCC_net_1, 
        F_AWADDR_HADDR0(4) => VCC_net_1, F_AWADDR_HADDR0(3) => 
        VCC_net_1, F_AWADDR_HADDR0(2) => VCC_net_1, 
        F_AWADDR_HADDR0(1) => VCC_net_1, F_AWADDR_HADDR0(0) => 
        VCC_net_1, F_AWBURST_HTRANS0(1) => GND_net_1, 
        F_AWBURST_HTRANS0(0) => GND_net_1, F_AWID_HSEL0(3) => 
        GND_net_1, F_AWID_HSEL0(2) => GND_net_1, F_AWID_HSEL0(1)
         => GND_net_1, F_AWID_HSEL0(0) => GND_net_1, 
        F_AWLEN_HBURST0(3) => GND_net_1, F_AWLEN_HBURST0(2) => 
        GND_net_1, F_AWLEN_HBURST0(1) => GND_net_1, 
        F_AWLEN_HBURST0(0) => GND_net_1, F_AWLOCK_HMASTLOCK0(1)
         => GND_net_1, F_AWLOCK_HMASTLOCK0(0) => GND_net_1, 
        F_AWSIZE_HSIZE0(1) => GND_net_1, F_AWSIZE_HSIZE0(0) => 
        GND_net_1, F_AWVALID_HWRITE0 => GND_net_1, F_BREADY => 
        GND_net_1, F_RMW_AXI => GND_net_1, F_RREADY => GND_net_1, 
        F_WDATA_HWDATA01(63) => VCC_net_1, F_WDATA_HWDATA01(62)
         => VCC_net_1, F_WDATA_HWDATA01(61) => VCC_net_1, 
        F_WDATA_HWDATA01(60) => VCC_net_1, F_WDATA_HWDATA01(59)
         => VCC_net_1, F_WDATA_HWDATA01(58) => VCC_net_1, 
        F_WDATA_HWDATA01(57) => VCC_net_1, F_WDATA_HWDATA01(56)
         => VCC_net_1, F_WDATA_HWDATA01(55) => VCC_net_1, 
        F_WDATA_HWDATA01(54) => VCC_net_1, F_WDATA_HWDATA01(53)
         => VCC_net_1, F_WDATA_HWDATA01(52) => VCC_net_1, 
        F_WDATA_HWDATA01(51) => VCC_net_1, F_WDATA_HWDATA01(50)
         => VCC_net_1, F_WDATA_HWDATA01(49) => VCC_net_1, 
        F_WDATA_HWDATA01(48) => VCC_net_1, F_WDATA_HWDATA01(47)
         => VCC_net_1, F_WDATA_HWDATA01(46) => VCC_net_1, 
        F_WDATA_HWDATA01(45) => VCC_net_1, F_WDATA_HWDATA01(44)
         => VCC_net_1, F_WDATA_HWDATA01(43) => VCC_net_1, 
        F_WDATA_HWDATA01(42) => VCC_net_1, F_WDATA_HWDATA01(41)
         => VCC_net_1, F_WDATA_HWDATA01(40) => VCC_net_1, 
        F_WDATA_HWDATA01(39) => VCC_net_1, F_WDATA_HWDATA01(38)
         => VCC_net_1, F_WDATA_HWDATA01(37) => VCC_net_1, 
        F_WDATA_HWDATA01(36) => VCC_net_1, F_WDATA_HWDATA01(35)
         => VCC_net_1, F_WDATA_HWDATA01(34) => VCC_net_1, 
        F_WDATA_HWDATA01(33) => VCC_net_1, F_WDATA_HWDATA01(32)
         => VCC_net_1, F_WDATA_HWDATA01(31) => VCC_net_1, 
        F_WDATA_HWDATA01(30) => VCC_net_1, F_WDATA_HWDATA01(29)
         => VCC_net_1, F_WDATA_HWDATA01(28) => VCC_net_1, 
        F_WDATA_HWDATA01(27) => VCC_net_1, F_WDATA_HWDATA01(26)
         => VCC_net_1, F_WDATA_HWDATA01(25) => VCC_net_1, 
        F_WDATA_HWDATA01(24) => VCC_net_1, F_WDATA_HWDATA01(23)
         => VCC_net_1, F_WDATA_HWDATA01(22) => VCC_net_1, 
        F_WDATA_HWDATA01(21) => VCC_net_1, F_WDATA_HWDATA01(20)
         => VCC_net_1, F_WDATA_HWDATA01(19) => VCC_net_1, 
        F_WDATA_HWDATA01(18) => VCC_net_1, F_WDATA_HWDATA01(17)
         => VCC_net_1, F_WDATA_HWDATA01(16) => VCC_net_1, 
        F_WDATA_HWDATA01(15) => VCC_net_1, F_WDATA_HWDATA01(14)
         => VCC_net_1, F_WDATA_HWDATA01(13) => VCC_net_1, 
        F_WDATA_HWDATA01(12) => VCC_net_1, F_WDATA_HWDATA01(11)
         => VCC_net_1, F_WDATA_HWDATA01(10) => VCC_net_1, 
        F_WDATA_HWDATA01(9) => VCC_net_1, F_WDATA_HWDATA01(8) => 
        VCC_net_1, F_WDATA_HWDATA01(7) => VCC_net_1, 
        F_WDATA_HWDATA01(6) => VCC_net_1, F_WDATA_HWDATA01(5) => 
        VCC_net_1, F_WDATA_HWDATA01(4) => VCC_net_1, 
        F_WDATA_HWDATA01(3) => VCC_net_1, F_WDATA_HWDATA01(2) => 
        VCC_net_1, F_WDATA_HWDATA01(1) => VCC_net_1, 
        F_WDATA_HWDATA01(0) => VCC_net_1, F_WID_HREADY01(3) => 
        GND_net_1, F_WID_HREADY01(2) => GND_net_1, 
        F_WID_HREADY01(1) => GND_net_1, F_WID_HREADY01(0) => 
        GND_net_1, F_WLAST => GND_net_1, F_WSTRB(7) => GND_net_1, 
        F_WSTRB(6) => GND_net_1, F_WSTRB(5) => GND_net_1, 
        F_WSTRB(4) => GND_net_1, F_WSTRB(3) => GND_net_1, 
        F_WSTRB(2) => GND_net_1, F_WSTRB(1) => GND_net_1, 
        F_WSTRB(0) => GND_net_1, F_WVALID => GND_net_1, 
        FPGA_MDDR_ARESET_N => VCC_net_1, MDDR_FABRIC_PADDR(10)
         => CORECONFIGP_0_MDDR_APBmslave_PADDR(10), 
        MDDR_FABRIC_PADDR(9) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(9), 
        MDDR_FABRIC_PADDR(8) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(8), 
        MDDR_FABRIC_PADDR(7) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(7), 
        MDDR_FABRIC_PADDR(6) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(6), 
        MDDR_FABRIC_PADDR(5) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(5), 
        MDDR_FABRIC_PADDR(4) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(4), 
        MDDR_FABRIC_PADDR(3) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(3), 
        MDDR_FABRIC_PADDR(2) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(2), 
        MDDR_FABRIC_PENABLE => 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE, MDDR_FABRIC_PSEL
         => CORECONFIGP_0_MDDR_APBmslave_PSELx, 
        MDDR_FABRIC_PWDATA(15) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(15), 
        MDDR_FABRIC_PWDATA(14) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(14), 
        MDDR_FABRIC_PWDATA(13) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(13), 
        MDDR_FABRIC_PWDATA(12) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(12), 
        MDDR_FABRIC_PWDATA(11) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(11), 
        MDDR_FABRIC_PWDATA(10) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(10), 
        MDDR_FABRIC_PWDATA(9) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(9), 
        MDDR_FABRIC_PWDATA(8) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(8), 
        MDDR_FABRIC_PWDATA(7) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(7), 
        MDDR_FABRIC_PWDATA(6) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(6), 
        MDDR_FABRIC_PWDATA(5) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(5), 
        MDDR_FABRIC_PWDATA(4) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(4), 
        MDDR_FABRIC_PWDATA(3) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(3), 
        MDDR_FABRIC_PWDATA(2) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(2), 
        MDDR_FABRIC_PWDATA(1) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(1), 
        MDDR_FABRIC_PWDATA(0) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(0), 
        MDDR_FABRIC_PWRITE => CORECONFIGP_0_MDDR_APBmslave_PWRITE, 
        PRESET_N => \CORECONFIGP_0_APB_S_PRESET_N\, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_IN => GPIO_GPIO_3_BI_PAD_Y, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN => GPIO_GPIO_4_BI_PAD_Y, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_IN => GND_net_1, DM_IN(2)
         => GND_net_1, DM_IN(1) => MDDR_DM_RDQS_1_PAD_Y, DM_IN(0)
         => MDDR_DM_RDQS_0_PAD_Y, DRAM_DQ_IN(17) => GND_net_1, 
        DRAM_DQ_IN(16) => GND_net_1, DRAM_DQ_IN(15) => 
        MDDR_DQ_15_PAD_Y, DRAM_DQ_IN(14) => MDDR_DQ_14_PAD_Y, 
        DRAM_DQ_IN(13) => MDDR_DQ_13_PAD_Y, DRAM_DQ_IN(12) => 
        MDDR_DQ_12_PAD_Y, DRAM_DQ_IN(11) => MDDR_DQ_11_PAD_Y, 
        DRAM_DQ_IN(10) => MDDR_DQ_10_PAD_Y, DRAM_DQ_IN(9) => 
        MDDR_DQ_9_PAD_Y, DRAM_DQ_IN(8) => MDDR_DQ_8_PAD_Y, 
        DRAM_DQ_IN(7) => MDDR_DQ_7_PAD_Y, DRAM_DQ_IN(6) => 
        MDDR_DQ_6_PAD_Y, DRAM_DQ_IN(5) => MDDR_DQ_5_PAD_Y, 
        DRAM_DQ_IN(4) => MDDR_DQ_4_PAD_Y, DRAM_DQ_IN(3) => 
        MDDR_DQ_3_PAD_Y, DRAM_DQ_IN(2) => MDDR_DQ_2_PAD_Y, 
        DRAM_DQ_IN(1) => MDDR_DQ_1_PAD_Y, DRAM_DQ_IN(0) => 
        MDDR_DQ_0_PAD_Y, DRAM_DQS_IN(2) => GND_net_1, 
        DRAM_DQS_IN(1) => MDDR_DQS_1_PAD_Y, DRAM_DQS_IN(0) => 
        MDDR_DQS_0_PAD_Y, DRAM_FIFO_WE_IN(1) => GND_net_1, 
        DRAM_FIFO_WE_IN(0) => MDDR_DQS_TMATCH_0_IN_PAD_Y, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_IN => GND_net_1, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_IN => GND_net_1, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_IN => I2C_1_SCL_PAD_Y, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_IN => I2C_1_SDA_PAD_Y, 
        MGPIO0B_IN => GPIO_GPIO_0_BI_PAD_Y, MGPIO10B_IN => 
        GND_net_1, MGPIO1B_IN => GND_net_1, MGPIO25A_IN => 
        GPIO_GPIO_25_BI_PAD_Y, MGPIO26A_IN => 
        GPIO_GPIO_26_BI_PAD_Y, MGPIO27A_IN => GND_net_1, 
        MGPIO28A_IN => GND_net_1, MGPIO29A_IN => GND_net_1, 
        MGPIO2B_IN => GND_net_1, MGPIO30A_IN => GND_net_1, 
        MGPIO31A_IN => GPIO_GPIO_31_BI_PAD_Y, MGPIO3B_IN => 
        GND_net_1, MGPIO4B_IN => GND_net_1, MGPIO5B_IN => 
        GND_net_1, MGPIO6B_IN => GND_net_1, MGPIO7B_IN => 
        GND_net_1, MGPIO8B_IN => GND_net_1, MGPIO9B_IN => 
        GND_net_1, MMUART0_CTS_USBC_DATA7_MGPIO19B_IN => 
        GND_net_1, MMUART0_DCD_MGPIO22B_IN => GND_net_1, 
        MMUART0_DSR_MGPIO20B_IN => GND_net_1, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_IN => GND_net_1, 
        MMUART0_RI_MGPIO21B_IN => GND_net_1, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_IN => GND_net_1, 
        MMUART0_RXD_USBC_STP_MGPIO28B_IN => GND_net_1, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_IN => GND_net_1, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_IN => GND_net_1, 
        MMUART1_CTS_MGPIO13B_IN => GND_net_1, 
        MMUART1_DCD_MGPIO16B_IN => GPIO_GPIO_16_BI_PAD_Y, 
        MMUART1_DSR_MGPIO14B_IN => GPIO_GPIO_14_BI_PAD_Y, 
        MMUART1_DTR_MGPIO12B_IN => GPIO_GPIO_12_BI_PAD_Y, 
        MMUART1_RI_MGPIO15B_IN => GPIO_GPIO_15_BI_PAD_Y, 
        MMUART1_RTS_MGPIO11B_IN => GND_net_1, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_IN => MMUART_1_RXD_PAD_Y, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_IN => GND_net_1, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_IN => GND_net_1, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN => GND_net_1, 
        RGMII_MDC_RMII_MDC_IN => GND_net_1, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN => GND_net_1, 
        RGMII_RX_CLK_IN => GND_net_1, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN => GND_net_1, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN => GND_net_1, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN => GND_net_1, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN => GND_net_1, 
        RGMII_RXD3_USBB_DATA4_IN => GND_net_1, RGMII_TX_CLK_IN
         => GND_net_1, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN => 
        GND_net_1, RGMII_TXD0_RMII_TXD0_USBB_DIR_IN => GND_net_1, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_IN => GND_net_1, 
        RGMII_TXD2_USBB_DATA5_IN => GND_net_1, 
        RGMII_TXD3_USBB_DATA6_IN => GND_net_1, 
        SPI0_SCK_USBA_XCLK_IN => SPI_0_CLK_PAD_Y, 
        SPI0_SDI_USBA_DIR_MGPIO5A_IN => SPI_0_DI_PAD_Y, 
        SPI0_SDO_USBA_STP_MGPIO6A_IN => GND_net_1, 
        SPI0_SS0_USBA_NXT_MGPIO7A_IN => SPI_0_SS0_PAD_Y, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_IN => GND_net_1, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_IN => GND_net_1, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_IN => GND_net_1, 
        SPI0_SS4_MGPIO19A_IN => GND_net_1, SPI0_SS5_MGPIO20A_IN
         => GND_net_1, SPI0_SS6_MGPIO21A_IN => GND_net_1, 
        SPI0_SS7_MGPIO22A_IN => GND_net_1, SPI1_SCK_IN => 
        GND_net_1, SPI1_SDI_MGPIO11A_IN => GND_net_1, 
        SPI1_SDO_MGPIO12A_IN => GND_net_1, SPI1_SS0_MGPIO13A_IN
         => GND_net_1, SPI1_SS1_MGPIO14A_IN => GND_net_1, 
        SPI1_SS2_MGPIO15A_IN => GND_net_1, SPI1_SS3_MGPIO16A_IN
         => GND_net_1, SPI1_SS4_MGPIO17A_IN => 
        GPIO_GPIO_17_BI_PAD_Y, SPI1_SS5_MGPIO18A_IN => 
        GPIO_GPIO_18_BI_PAD_Y, SPI1_SS6_MGPIO23A_IN => GND_net_1, 
        SPI1_SS7_MGPIO24A_IN => GND_net_1, USBC_XCLK_IN => 
        GND_net_1, USBD_DATA0_IN => GND_net_1, USBD_DATA1_IN => 
        GND_net_1, USBD_DATA2_IN => GND_net_1, USBD_DATA3_IN => 
        GND_net_1, USBD_DATA4_IN => GND_net_1, USBD_DATA5_IN => 
        GND_net_1, USBD_DATA6_IN => GND_net_1, 
        USBD_DATA7_MGPIO23B_IN => GND_net_1, USBD_DIR_IN => 
        GND_net_1, USBD_NXT_IN => GND_net_1, USBD_STP_IN => 
        GND_net_1, USBD_XCLK_IN => GND_net_1, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT => 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT => 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT => OPEN, DRAM_ADDR(15)
         => \DRAM_ADDR_net_0[15]\, DRAM_ADDR(14) => 
        \DRAM_ADDR_net_0[14]\, DRAM_ADDR(13) => 
        \DRAM_ADDR_net_0[13]\, DRAM_ADDR(12) => 
        \DRAM_ADDR_net_0[12]\, DRAM_ADDR(11) => 
        \DRAM_ADDR_net_0[11]\, DRAM_ADDR(10) => 
        \DRAM_ADDR_net_0[10]\, DRAM_ADDR(9) => 
        \DRAM_ADDR_net_0[9]\, DRAM_ADDR(8) => 
        \DRAM_ADDR_net_0[8]\, DRAM_ADDR(7) => 
        \DRAM_ADDR_net_0[7]\, DRAM_ADDR(6) => 
        \DRAM_ADDR_net_0[6]\, DRAM_ADDR(5) => 
        \DRAM_ADDR_net_0[5]\, DRAM_ADDR(4) => 
        \DRAM_ADDR_net_0[4]\, DRAM_ADDR(3) => 
        \DRAM_ADDR_net_0[3]\, DRAM_ADDR(2) => 
        \DRAM_ADDR_net_0[2]\, DRAM_ADDR(1) => 
        \DRAM_ADDR_net_0[1]\, DRAM_ADDR(0) => 
        \DRAM_ADDR_net_0[0]\, DRAM_BA(2) => \DRAM_BA_net_0[2]\, 
        DRAM_BA(1) => \DRAM_BA_net_0[1]\, DRAM_BA(0) => 
        \DRAM_BA_net_0[0]\, DRAM_CASN => MSS_ADLIB_INST_DRAM_CASN, 
        DRAM_CKE => MSS_ADLIB_INST_DRAM_CKE, DRAM_CLK => 
        MSS_ADLIB_INST_DRAM_CLK, DRAM_CSN => 
        MSS_ADLIB_INST_DRAM_CSN, DRAM_DM_RDQS_OUT(2) => nc22, 
        DRAM_DM_RDQS_OUT(1) => \DRAM_DM_RDQS_OUT_net_0[1]\, 
        DRAM_DM_RDQS_OUT(0) => \DRAM_DM_RDQS_OUT_net_0[0]\, 
        DRAM_DQ_OUT(17) => nc210, DRAM_DQ_OUT(16) => nc185, 
        DRAM_DQ_OUT(15) => \DRAM_DQ_OUT_net_0[15]\, 
        DRAM_DQ_OUT(14) => \DRAM_DQ_OUT_net_0[14]\, 
        DRAM_DQ_OUT(13) => \DRAM_DQ_OUT_net_0[13]\, 
        DRAM_DQ_OUT(12) => \DRAM_DQ_OUT_net_0[12]\, 
        DRAM_DQ_OUT(11) => \DRAM_DQ_OUT_net_0[11]\, 
        DRAM_DQ_OUT(10) => \DRAM_DQ_OUT_net_0[10]\, 
        DRAM_DQ_OUT(9) => \DRAM_DQ_OUT_net_0[9]\, DRAM_DQ_OUT(8)
         => \DRAM_DQ_OUT_net_0[8]\, DRAM_DQ_OUT(7) => 
        \DRAM_DQ_OUT_net_0[7]\, DRAM_DQ_OUT(6) => 
        \DRAM_DQ_OUT_net_0[6]\, DRAM_DQ_OUT(5) => 
        \DRAM_DQ_OUT_net_0[5]\, DRAM_DQ_OUT(4) => 
        \DRAM_DQ_OUT_net_0[4]\, DRAM_DQ_OUT(3) => 
        \DRAM_DQ_OUT_net_0[3]\, DRAM_DQ_OUT(2) => 
        \DRAM_DQ_OUT_net_0[2]\, DRAM_DQ_OUT(1) => 
        \DRAM_DQ_OUT_net_0[1]\, DRAM_DQ_OUT(0) => 
        \DRAM_DQ_OUT_net_0[0]\, DRAM_DQS_OUT(2) => nc143, 
        DRAM_DQS_OUT(1) => \DRAM_DQS_OUT_net_0[1]\, 
        DRAM_DQS_OUT(0) => \DRAM_DQS_OUT_net_0[0]\, 
        DRAM_FIFO_WE_OUT(1) => nc77, DRAM_FIFO_WE_OUT(0) => 
        \DRAM_FIFO_WE_OUT_net_0[0]\, DRAM_ODT => 
        MSS_ADLIB_INST_DRAM_ODT, DRAM_RASN => 
        MSS_ADLIB_INST_DRAM_RASN, DRAM_RSTN => 
        MSS_ADLIB_INST_DRAM_RSTN, DRAM_WEN => 
        MSS_ADLIB_INST_DRAM_WEN, I2C0_SCL_USBC_DATA1_MGPIO31B_OUT
         => OPEN, I2C0_SDA_USBC_DATA0_MGPIO30B_OUT => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OUT => 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OUT => 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT, 
        MGPIO0B_OUT => MSS_ADLIB_INST_MGPIO0B_OUT, MGPIO10B_OUT
         => OPEN, MGPIO1B_OUT => OPEN, MGPIO25A_OUT => 
        MSS_ADLIB_INST_MGPIO25A_OUT, MGPIO26A_OUT => 
        MSS_ADLIB_INST_MGPIO26A_OUT, MGPIO27A_OUT => OPEN, 
        MGPIO28A_OUT => OPEN, MGPIO29A_OUT => OPEN, MGPIO2B_OUT
         => OPEN, MGPIO30A_OUT => OPEN, MGPIO31A_OUT => 
        MSS_ADLIB_INST_MGPIO31A_OUT, MGPIO3B_OUT => OPEN, 
        MGPIO4B_OUT => OPEN, MGPIO5B_OUT => OPEN, MGPIO6B_OUT => 
        OPEN, MGPIO7B_OUT => OPEN, MGPIO8B_OUT => OPEN, 
        MGPIO9B_OUT => OPEN, MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT
         => OPEN, MMUART0_DCD_MGPIO22B_OUT => OPEN, 
        MMUART0_DSR_MGPIO20B_OUT => OPEN, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT => OPEN, 
        MMUART0_RI_MGPIO21B_OUT => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OUT => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OUT => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OUT => OPEN, 
        MMUART1_CTS_MGPIO13B_OUT => OPEN, 
        MMUART1_DCD_MGPIO16B_OUT => 
        MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OUT, 
        MMUART1_DSR_MGPIO14B_OUT => 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OUT, 
        MMUART1_DTR_MGPIO12B_OUT => 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OUT, 
        MMUART1_RI_MGPIO15B_OUT => 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OUT, 
        MMUART1_RTS_MGPIO11B_OUT => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT => OPEN, 
        RGMII_MDC_RMII_MDC_OUT => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT => OPEN, 
        RGMII_RX_CLK_OUT => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT => OPEN, 
        RGMII_RXD3_USBB_DATA4_OUT => OPEN, RGMII_TX_CLK_OUT => 
        OPEN, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OUT => OPEN, 
        RGMII_TXD2_USBB_DATA5_OUT => OPEN, 
        RGMII_TXD3_USBB_DATA6_OUT => OPEN, SPI0_SCK_USBA_XCLK_OUT
         => MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, 
        SPI0_SDI_USBA_DIR_MGPIO5A_OUT => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OUT => 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OUT => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OUT => 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OUT, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OUT => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OUT => OPEN, 
        SPI0_SS4_MGPIO19A_OUT => OPEN, SPI0_SS5_MGPIO20A_OUT => 
        MSS_ADLIB_INST_SPI0_SS5_MGPIO20A_OUT, 
        SPI0_SS6_MGPIO21A_OUT => OPEN, SPI0_SS7_MGPIO22A_OUT => 
        OPEN, SPI1_SCK_OUT => OPEN, SPI1_SDI_MGPIO11A_OUT => OPEN, 
        SPI1_SDO_MGPIO12A_OUT => OPEN, SPI1_SS0_MGPIO13A_OUT => 
        OPEN, SPI1_SS1_MGPIO14A_OUT => OPEN, 
        SPI1_SS2_MGPIO15A_OUT => OPEN, SPI1_SS3_MGPIO16A_OUT => 
        OPEN, SPI1_SS4_MGPIO17A_OUT => 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OUT, 
        SPI1_SS5_MGPIO18A_OUT => 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OUT, 
        SPI1_SS6_MGPIO23A_OUT => OPEN, SPI1_SS7_MGPIO24A_OUT => 
        OPEN, USBC_XCLK_OUT => OPEN, USBD_DATA0_OUT => OPEN, 
        USBD_DATA1_OUT => OPEN, USBD_DATA2_OUT => OPEN, 
        USBD_DATA3_OUT => OPEN, USBD_DATA4_OUT => OPEN, 
        USBD_DATA5_OUT => OPEN, USBD_DATA6_OUT => OPEN, 
        USBD_DATA7_MGPIO23B_OUT => OPEN, USBD_DIR_OUT => OPEN, 
        USBD_NXT_OUT => OPEN, USBD_STP_OUT => OPEN, USBD_XCLK_OUT
         => OPEN, CAN_RXBUS_USBA_DATA1_MGPIO3A_OE => 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OE, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE => 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OE => OPEN, DM_OE(2) => nc6, 
        DM_OE(1) => \DM_OE_net_0[1]\, DM_OE(0) => 
        \DM_OE_net_0[0]\, DRAM_DQ_OE(17) => nc109, DRAM_DQ_OE(16)
         => nc87, DRAM_DQ_OE(15) => \DRAM_DQ_OE_net_0[15]\, 
        DRAM_DQ_OE(14) => \DRAM_DQ_OE_net_0[14]\, DRAM_DQ_OE(13)
         => \DRAM_DQ_OE_net_0[13]\, DRAM_DQ_OE(12) => 
        \DRAM_DQ_OE_net_0[12]\, DRAM_DQ_OE(11) => 
        \DRAM_DQ_OE_net_0[11]\, DRAM_DQ_OE(10) => 
        \DRAM_DQ_OE_net_0[10]\, DRAM_DQ_OE(9) => 
        \DRAM_DQ_OE_net_0[9]\, DRAM_DQ_OE(8) => 
        \DRAM_DQ_OE_net_0[8]\, DRAM_DQ_OE(7) => 
        \DRAM_DQ_OE_net_0[7]\, DRAM_DQ_OE(6) => 
        \DRAM_DQ_OE_net_0[6]\, DRAM_DQ_OE(5) => 
        \DRAM_DQ_OE_net_0[5]\, DRAM_DQ_OE(4) => 
        \DRAM_DQ_OE_net_0[4]\, DRAM_DQ_OE(3) => 
        \DRAM_DQ_OE_net_0[3]\, DRAM_DQ_OE(2) => 
        \DRAM_DQ_OE_net_0[2]\, DRAM_DQ_OE(1) => 
        \DRAM_DQ_OE_net_0[1]\, DRAM_DQ_OE(0) => 
        \DRAM_DQ_OE_net_0[0]\, DRAM_DQS_OE(2) => nc123, 
        DRAM_DQS_OE(1) => \DRAM_DQS_OE_net_0[1]\, DRAM_DQS_OE(0)
         => \DRAM_DQS_OE_net_0[0]\, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_OE => OPEN, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OE => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OE => 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OE => 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE, MGPIO0B_OE
         => MSS_ADLIB_INST_MGPIO0B_OE, MGPIO10B_OE => OPEN, 
        MGPIO1B_OE => OPEN, MGPIO25A_OE => 
        MSS_ADLIB_INST_MGPIO25A_OE, MGPIO26A_OE => 
        MSS_ADLIB_INST_MGPIO26A_OE, MGPIO27A_OE => OPEN, 
        MGPIO28A_OE => OPEN, MGPIO29A_OE => OPEN, MGPIO2B_OE => 
        OPEN, MGPIO30A_OE => OPEN, MGPIO31A_OE => 
        MSS_ADLIB_INST_MGPIO31A_OE, MGPIO3B_OE => OPEN, 
        MGPIO4B_OE => OPEN, MGPIO5B_OE => OPEN, MGPIO6B_OE => 
        OPEN, MGPIO7B_OE => OPEN, MGPIO8B_OE => OPEN, MGPIO9B_OE
         => OPEN, MMUART0_CTS_USBC_DATA7_MGPIO19B_OE => OPEN, 
        MMUART0_DCD_MGPIO22B_OE => OPEN, MMUART0_DSR_MGPIO20B_OE
         => OPEN, MMUART0_DTR_USBC_DATA6_MGPIO18B_OE => OPEN, 
        MMUART0_RI_MGPIO21B_OE => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OE => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OE => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OE => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OE => OPEN, 
        MMUART1_CTS_MGPIO13B_OE => OPEN, MMUART1_DCD_MGPIO16B_OE
         => MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OE, 
        MMUART1_DSR_MGPIO14B_OE => 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OE, 
        MMUART1_DTR_MGPIO12B_OE => 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OE, 
        MMUART1_RI_MGPIO15B_OE => 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OE, 
        MMUART1_RTS_MGPIO11B_OE => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OE => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OE => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OE => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE => OPEN, 
        RGMII_MDC_RMII_MDC_OE => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE => OPEN, 
        RGMII_RX_CLK_OE => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE => OPEN, 
        RGMII_RXD3_USBB_DATA4_OE => OPEN, RGMII_TX_CLK_OE => OPEN, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OE => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OE => OPEN, 
        RGMII_TXD2_USBB_DATA5_OE => OPEN, 
        RGMII_TXD3_USBB_DATA6_OE => OPEN, SPI0_SCK_USBA_XCLK_OE
         => MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, 
        SPI0_SDI_USBA_DIR_MGPIO5A_OE => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OE => 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OE => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OE => 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OE, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OE => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OE => OPEN, 
        SPI0_SS4_MGPIO19A_OE => OPEN, SPI0_SS5_MGPIO20A_OE => 
        OPEN, SPI0_SS6_MGPIO21A_OE => OPEN, SPI0_SS7_MGPIO22A_OE
         => OPEN, SPI1_SCK_OE => OPEN, SPI1_SDI_MGPIO11A_OE => 
        OPEN, SPI1_SDO_MGPIO12A_OE => OPEN, SPI1_SS0_MGPIO13A_OE
         => OPEN, SPI1_SS1_MGPIO14A_OE => OPEN, 
        SPI1_SS2_MGPIO15A_OE => OPEN, SPI1_SS3_MGPIO16A_OE => 
        OPEN, SPI1_SS4_MGPIO17A_OE => 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OE, SPI1_SS5_MGPIO18A_OE
         => MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OE, 
        SPI1_SS6_MGPIO23A_OE => OPEN, SPI1_SS7_MGPIO24A_OE => 
        OPEN, USBC_XCLK_OE => OPEN, USBD_DATA0_OE => OPEN, 
        USBD_DATA1_OE => OPEN, USBD_DATA2_OE => OPEN, 
        USBD_DATA3_OE => OPEN, USBD_DATA4_OE => OPEN, 
        USBD_DATA5_OE => OPEN, USBD_DATA6_OE => OPEN, 
        USBD_DATA7_MGPIO23B_OE => OPEN, USBD_DIR_OE => OPEN, 
        USBD_NXT_OE => OPEN, USBD_STP_OE => OPEN, USBD_XCLK_OE
         => OPEN);
    
    MDDR_RAS_N_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_RASN, PAD => MDDR_RAS_N);
    
    SPI_0_CLK_PAD : BIBUF
      port map(PAD => SPI_0_CLK, D => 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, E => 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, Y => 
        SPI_0_CLK_PAD_Y);
    
    MDDR_DQ_4_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(4), D => \DRAM_DQ_OUT_net_0[4]\, E
         => \DRAM_DQ_OE_net_0[4]\, Y => MDDR_DQ_4_PAD_Y);
    
    GPIO_GPIO_18_BI_PAD : BIBUF
      port map(PAD => GPIO_18_BI, D => 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OUT, E => 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OE, Y => 
        GPIO_GPIO_18_BI_PAD_Y);
    
    GPIO_GPIO_16_BI_PAD : BIBUF
      port map(PAD => GPIO_16_BI, D => 
        MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OE, Y => 
        GPIO_GPIO_16_BI_PAD_Y);
    
    MDDR_ADDR_10_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[10]\, PAD => MDDR_ADDR(10));
    
    MDDR_DQS_TMATCH_0_IN_PAD : INBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQS_TMATCH_0_IN, Y => 
        MDDR_DQS_TMATCH_0_IN_PAD_Y);
    
    MDDR_CS_N_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_CSN, PAD => MDDR_CS_N);
    
    MDDR_ADDR_4_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[4]\, PAD => MDDR_ADDR(4));
    
    SPI_0_SS0_PAD : BIBUF
      port map(PAD => SPI_0_SS0, D => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, E => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, Y => 
        SPI_0_SS0_PAD_Y);
    
    MDDR_DQ_7_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(7), D => \DRAM_DQ_OUT_net_0[7]\, E
         => \DRAM_DQ_OE_net_0[7]\, Y => MDDR_DQ_7_PAD_Y);
    
    MDDR_WE_N_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_WEN, PAD => MDDR_WE_N);
    
    MDDR_ADDR_8_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[8]\, PAD => MDDR_ADDR(8));
    
    GPIO_GPIO_3_BI_PAD : BIBUF
      port map(PAD => GPIO_3_BI, D => 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT, E => 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OE, Y => 
        GPIO_GPIO_3_BI_PAD_Y);
    
    MDDR_ADDR_15_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[15]\, PAD => MDDR_ADDR(15));
    
    MDDR_ADDR_0_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[0]\, PAD => MDDR_ADDR(0));
    
    MDDR_ADDR_1_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[1]\, PAD => MDDR_ADDR(1));
    
    GPIO_GPIO_20_OUT_PAD : OUTBUF
      port map(D => MSS_ADLIB_INST_SPI0_SS5_MGPIO20A_OUT, PAD => 
        GPIO_20_OUT);
    
    SPI_0_SS1_PAD : TRIBUFF
      port map(D => 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OUT, E => 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OE, PAD => 
        SPI_0_SS1);
    
    FIC_2_APB_M_PCLK_inferred_clock_RNIPG5 : CLKINT
      port map(A => FIC_2_APB_M_PCLK, Y => 
        \CORECONFIGP_0_APB_S_PCLK\);
    
    MDDR_DQ_13_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(13), D => \DRAM_DQ_OUT_net_0[13]\, 
        E => \DRAM_DQ_OE_net_0[13]\, Y => MDDR_DQ_13_PAD_Y);
    
    MDDR_ADDR_3_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[3]\, PAD => MDDR_ADDR(3));
    
    MMUART_1_RXD_PAD : INBUF
      port map(PAD => MMUART_1_RXD, Y => MMUART_1_RXD_PAD_Y);
    
    MDDR_BA_0_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_BA_net_0[0]\, PAD => MDDR_BA(0));
    
    GPIO_GPIO_26_BI_PAD : BIBUF
      port map(PAD => GPIO_26_BI, D => 
        MSS_ADLIB_INST_MGPIO26A_OUT, E => 
        MSS_ADLIB_INST_MGPIO26A_OE, Y => GPIO_GPIO_26_BI_PAD_Y);
    
    MDDR_DQ_6_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(6), D => \DRAM_DQ_OUT_net_0[6]\, E
         => \DRAM_DQ_OE_net_0[6]\, Y => MDDR_DQ_6_PAD_Y);
    
    MDDR_CLK_PAD : OUTBUF_DIFF
      generic map(IOSTD => "LPDDRI")

      port map(D => MSS_ADLIB_INST_DRAM_CLK, PADP => MDDR_CLK, 
        PADN => MDDR_CLK_N);
    
    MDDR_DQ_14_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(14), D => \DRAM_DQ_OUT_net_0[14]\, 
        E => \DRAM_DQ_OE_net_0[14]\, Y => MDDR_DQ_14_PAD_Y);
    
    GPIO_GPIO_15_BI_PAD : BIBUF
      port map(PAD => GPIO_15_BI, D => 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OE, Y => 
        GPIO_GPIO_15_BI_PAD_Y);
    
    MDDR_DQS_TMATCH_0_OUT_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_FIFO_WE_OUT_net_0[0]\, PAD => 
        MDDR_DQS_TMATCH_0_OUT);
    
    MDDR_BA_1_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_BA_net_0[1]\, PAD => MDDR_BA(1));
    
    MDDR_DQ_5_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(5), D => \DRAM_DQ_OUT_net_0[5]\, E
         => \DRAM_DQ_OE_net_0[5]\, Y => MDDR_DQ_5_PAD_Y);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreResetP is

    port( CORECONFIGP_0_CONFIG2_DONE              : in    std_logic;
          CORECONFIGP_0_CONFIG1_DONE              : in    std_logic;
          CORECONFIGP_0_APB_S_PRESET_N            : in    std_logic;
          m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F : in    std_logic;
          m2s010_som_sb_0_POWER_ON_RESET_N        : in    std_logic;
          INIT_DONE                               : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_O2F             : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz               : in    std_logic
        );

end CoreResetP;

architecture DEF_ARCH of CoreResetP is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \sm0_areset_n_rcosc\, sm0_areset_n_rcosc_0, 
        \sm0_areset_n_clk_base\, sm0_areset_n_clk_base_0, 
        \count_ddr[0]_net_1\, \count_ddr_s[0]\, \mss_ready_state\, 
        VCC_net_1, \POWER_ON_RESET_N_clk_base\, 
        \RESET_N_M2F_clk_base\, GND_net_1, \ddr_settled\, 
        \un14_count_ddr\, \count_ddr_enable\, 
        next_count_ddr_enable_0_sqmuxa, 
        \un1_next_ddr_ready_0_sqmuxa\, \mss_ready_select\, 
        \un6_fic_2_apb_m_preset_n_clk_base\, \sm0_state[0]_net_1\, 
        \sm0_state[6]_net_1\, \sm0_state[5]_net_1\, 
        \sm0_state[4]_net_1\, \sm0_state_ns[2]_net_1\, 
        \sm0_state[3]_net_1\, \sm0_state_ns[3]_net_1\, 
        \sm0_state[2]_net_1\, \sm0_state_ns[4]_net_1\, 
        \sm0_state[1]_net_1\, \sm0_state_ns[5]_net_1\, 
        \sm0_state_ns_a3[6]_net_1\, \MSS_HPMS_READY_int\, 
        \MSS_HPMS_READY_int_3\, sm0_areset_n_rcosc_q1, 
        sm0_areset_n_i_i, \release_sdif0_core_q1\, 
        \release_sdif0_core\, \POWER_ON_RESET_N_q1\, 
        \RESET_N_M2F_q1\, \FIC_2_APB_M_PRESET_N_q1\, 
        \sdif3_spll_lock_q1\, \count_ddr_enable_rcosc\, 
        \count_ddr_enable_q1\, \ddr_settled_clk_base\, 
        \ddr_settled_q1\, \release_sdif0_core_clk_base\, 
        \FIC_2_APB_M_PRESET_N_clk_base\, \sm0_areset_n_q1\, 
        \CONFIG1_DONE_clk_base\, \CONFIG1_DONE_q1\, 
        \CONFIG2_DONE_clk_base\, \CONFIG2_DONE_q1\, 
        \sdif3_spll_lock_q2\, \count_ddr[1]_net_1\, 
        \count_ddr_s[1]\, \count_ddr[2]_net_1\, \count_ddr_s[2]\, 
        \count_ddr[3]_net_1\, \count_ddr_s[3]\, 
        \count_ddr[4]_net_1\, \count_ddr_s[4]\, 
        \count_ddr[5]_net_1\, \count_ddr_s[5]\, 
        \count_ddr[6]_net_1\, \count_ddr_s[6]\, 
        \count_ddr[7]_net_1\, \count_ddr_s[7]\, 
        \count_ddr[8]_net_1\, \count_ddr_s[8]\, 
        \count_ddr[9]_net_1\, \count_ddr_s[9]\, 
        \count_ddr[10]_net_1\, \count_ddr_s[10]\, 
        \count_ddr[11]_net_1\, \count_ddr_s[11]\, 
        \count_ddr[12]_net_1\, \count_ddr_s[12]\, 
        \count_ddr[13]_net_1\, \count_ddr_s[13]_net_1\, 
        count_ddr_s_265_FCO, \count_ddr_cry[1]_net_1\, 
        \count_ddr_cry[2]_net_1\, \count_ddr_cry[3]_net_1\, 
        \count_ddr_cry[4]_net_1\, \count_ddr_cry[5]_net_1\, 
        \count_ddr_cry[6]_net_1\, \count_ddr_cry[7]_net_1\, 
        \count_ddr_cry[8]_net_1\, \count_ddr_cry[9]_net_1\, 
        \count_ddr_cry[10]_net_1\, \count_ddr_cry[11]_net_1\, 
        \count_ddr_cry[12]_net_1\, \un14_count_ddr_6\, 
        \un8_ddr_settled_clk_base\, \un14_count_ddr_9\, 
        \un14_count_ddr_8\, \un14_count_ddr_7\ : std_logic;

begin 


    un14_count_ddr : CFG4
      generic map(INIT => x"8000")

      port map(A => \un14_count_ddr_7\, B => \un14_count_ddr_6\, 
        C => \un14_count_ddr_8\, D => \un14_count_ddr_9\, Y => 
        \un14_count_ddr\);
    
    \sm0_state_ns[4]\ : CFG4
      generic map(INIT => x"FF70")

      port map(A => \release_sdif0_core_clk_base\, B => 
        \ddr_settled_clk_base\, C => \sm0_state[2]_net_1\, D => 
        next_count_ddr_enable_0_sqmuxa, Y => 
        \sm0_state_ns[4]_net_1\);
    
    sm0_areset_n_rcosc : SLE
      port map(D => sm0_areset_n_rcosc_q1, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => VCC_net_1, ALn => 
        sm0_areset_n_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        sm0_areset_n_rcosc_0);
    
    \count_ddr[3]\ : SLE
      port map(D => \count_ddr_s[3]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[3]_net_1\);
    
    sm0_areset_n_q1 : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => sm0_areset_n_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sm0_areset_n_q1\);
    
    MSS_HPMS_READY_int_RNINOKG : CFG2
      generic map(INIT => x"8")

      port map(A => \MSS_HPMS_READY_int\, B => 
        m2s010_som_sb_0_POWER_ON_RESET_N, Y => sm0_areset_n_i_i);
    
    count_ddr_enable_q1 : SLE
      port map(D => \count_ddr_enable\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => VCC_net_1, ALn => 
        \sm0_areset_n_rcosc\, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \count_ddr_enable_q1\);
    
    \sm0_state[6]\ : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => \sm0_areset_n_clk_base\, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sm0_state[6]_net_1\);
    
    \sm0_state[2]\ : SLE
      port map(D => \sm0_state_ns[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[2]_net_1\);
    
    FIC_2_APB_M_PRESET_N_clk_base : SLE
      port map(D => \FIC_2_APB_M_PRESET_N_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \FIC_2_APB_M_PRESET_N_clk_base\);
    
    \count_ddr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[3]_net_1\, S => \count_ddr_s[4]\, Y => 
        OPEN, FCO => \count_ddr_cry[4]_net_1\);
    
    un8_ddr_settled_clk_base : CFG2
      generic map(INIT => x"8")

      port map(A => \ddr_settled_clk_base\, B => 
        \release_sdif0_core_clk_base\, Y => 
        \un8_ddr_settled_clk_base\);
    
    INIT_DONE_int : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \sm0_state[0]_net_1\, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        INIT_DONE);
    
    \count_ddr[9]\ : SLE
      port map(D => \count_ddr_s[9]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[9]_net_1\);
    
    MSS_HPMS_READY_int : SLE
      port map(D => \MSS_HPMS_READY_int_3\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \MSS_HPMS_READY_int\);
    
    count_ddr_enable_rcosc : SLE
      port map(D => \count_ddr_enable_q1\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => VCC_net_1, ALn => 
        \sm0_areset_n_rcosc\, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \count_ddr_enable_rcosc\);
    
    sm0_areset_n_clk_base_RNIEFM9 : CLKINT
      port map(A => sm0_areset_n_clk_base_0, Y => 
        \sm0_areset_n_clk_base\);
    
    \count_ddr[7]\ : SLE
      port map(D => \count_ddr_s[7]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[7]_net_1\);
    
    \sm0_state_ns_a3[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \CONFIG2_DONE_clk_base\, B => 
        \sm0_state[1]_net_1\, Y => \sm0_state_ns_a3[6]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sm0_state[4]\ : SLE
      port map(D => \sm0_state_ns[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[4]_net_1\);
    
    MSS_HPMS_READY_int_3 : CFG3
      generic map(INIT => x"E0")

      port map(A => \RESET_N_M2F_clk_base\, B => 
        \mss_ready_select\, C => \FIC_2_APB_M_PRESET_N_clk_base\, 
        Y => \MSS_HPMS_READY_int_3\);
    
    count_ddr_enable : SLE
      port map(D => next_count_ddr_enable_0_sqmuxa, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        \un1_next_ddr_ready_0_sqmuxa\, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \count_ddr_enable\);
    
    \count_ddr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[9]_net_1\, S => \count_ddr_s[10]\, Y => 
        OPEN, FCO => \count_ddr_cry[10]_net_1\);
    
    \sm0_state[5]\ : SLE
      port map(D => \sm0_state[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[5]_net_1\);
    
    \count_ddr_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[10]_net_1\, S => \count_ddr_s[11]\, Y => 
        OPEN, FCO => \count_ddr_cry[11]_net_1\);
    
    \count_ddr[8]\ : SLE
      port map(D => \count_ddr_s[8]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[8]_net_1\);
    
    \sm0_state_ns[2]\ : CFG3
      generic map(INIT => x"AE")

      port map(A => \sm0_state[5]_net_1\, B => 
        \sm0_state[4]_net_1\, C => \CONFIG1_DONE_clk_base\, Y => 
        \sm0_state_ns[2]_net_1\);
    
    sm0_areset_n_clk_base : SLE
      port map(D => \sm0_areset_n_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        sm0_areset_n_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        sm0_areset_n_clk_base_0);
    
    \count_ddr_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[11]_net_1\, S => \count_ddr_s[12]\, Y => 
        OPEN, FCO => \count_ddr_cry[12]_net_1\);
    
    mss_ready_state : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \RESET_N_M2F_clk_base\, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_state\);
    
    \sm0_state[1]\ : SLE
      port map(D => \sm0_state_ns[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[1]_net_1\);
    
    next_count_ddr_enable_0_sqmuxa_0_a3 : CFG2
      generic map(INIT => x"8")

      port map(A => \sdif3_spll_lock_q2\, B => 
        \sm0_state[3]_net_1\, Y => next_count_ddr_enable_0_sqmuxa);
    
    ddr_settled_clk_base : SLE
      port map(D => \ddr_settled_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ddr_settled_clk_base\);
    
    FIC_2_APB_M_PRESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \FIC_2_APB_M_PRESET_N_q1\);
    
    un14_count_ddr_7 : CFG4
      generic map(INIT => x"8000")

      port map(A => \count_ddr[10]_net_1\, B => 
        \count_ddr[9]_net_1\, C => \count_ddr[8]_net_1\, D => 
        \count_ddr[4]_net_1\, Y => \un14_count_ddr_7\);
    
    \count_ddr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[7]_net_1\, S => \count_ddr_s[8]\, Y => 
        OPEN, FCO => \count_ddr_cry[8]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \count_ddr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \count_ddr[0]_net_1\, Y => \count_ddr_s[0]\);
    
    count_ddr_s_265 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => count_ddr_s_265_FCO);
    
    POWER_ON_RESET_N_clk_base : SLE
      port map(D => \POWER_ON_RESET_N_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        m2s010_som_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \POWER_ON_RESET_N_clk_base\);
    
    \count_ddr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => count_ddr_s_265_FCO, S
         => \count_ddr_s[1]\, Y => OPEN, FCO => 
        \count_ddr_cry[1]_net_1\);
    
    RESET_N_M2F_q1 : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RESET_N_M2F_q1\);
    
    release_sdif0_core_q1 : SLE
      port map(D => \release_sdif0_core\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \release_sdif0_core_q1\);
    
    \count_ddr[10]\ : SLE
      port map(D => \count_ddr_s[10]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[10]_net_1\);
    
    \count_ddr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[5]_net_1\, S => \count_ddr_s[6]\, Y => 
        OPEN, FCO => \count_ddr_cry[6]_net_1\);
    
    \count_ddr_s[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[12]_net_1\, S => \count_ddr_s[13]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \count_ddr[5]\ : SLE
      port map(D => \count_ddr_s[5]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[5]_net_1\);
    
    \count_ddr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[2]_net_1\, S => \count_ddr_s[3]\, Y => 
        OPEN, FCO => \count_ddr_cry[3]_net_1\);
    
    \count_ddr[2]\ : SLE
      port map(D => \count_ddr_s[2]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[2]_net_1\);
    
    sdif0_areset_n_rcosc_q1 : SLE
      port map(D => VCC_net_1, CLK => FABOSC_0_RCOSC_25_50MHZ_O2F, 
        EN => VCC_net_1, ALn => sm0_areset_n_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => sm0_areset_n_rcosc_q1);
    
    \count_ddr[1]\ : SLE
      port map(D => \count_ddr_s[1]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[1]_net_1\);
    
    \sm0_state[0]\ : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \sm0_state_ns_a3[6]_net_1\, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[0]_net_1\);
    
    un14_count_ddr_8 : CFG4
      generic map(INIT => x"0002")

      port map(A => \count_ddr[13]_net_1\, B => 
        \count_ddr[2]_net_1\, C => \count_ddr[1]_net_1\, D => 
        \count_ddr[0]_net_1\, Y => \un14_count_ddr_8\);
    
    \count_ddr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[1]_net_1\, S => \count_ddr_s[2]\, Y => 
        OPEN, FCO => \count_ddr_cry[2]_net_1\);
    
    \count_ddr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[4]_net_1\, S => \count_ddr_s[5]\, Y => 
        OPEN, FCO => \count_ddr_cry[5]_net_1\);
    
    ddr_settled_q1 : SLE
      port map(D => \ddr_settled\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ddr_settled_q1\);
    
    \count_ddr[11]\ : SLE
      port map(D => \count_ddr_s[11]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[11]_net_1\);
    
    un14_count_ddr_9 : CFG4
      generic map(INIT => x"0001")

      port map(A => \count_ddr[12]_net_1\, B => 
        \count_ddr[11]_net_1\, C => \count_ddr[5]_net_1\, D => 
        \count_ddr[3]_net_1\, Y => \un14_count_ddr_9\);
    
    \sm0_state[3]\ : SLE
      port map(D => \sm0_state_ns[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[3]_net_1\);
    
    \sm0_state_ns[3]\ : CFG4
      generic map(INIT => x"F222")

      port map(A => \sm0_state[3]_net_1\, B => 
        \sdif3_spll_lock_q2\, C => \sm0_state[4]_net_1\, D => 
        \CONFIG1_DONE_clk_base\, Y => \sm0_state_ns[3]_net_1\);
    
    \count_ddr[0]\ : SLE
      port map(D => \count_ddr_s[0]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[0]_net_1\);
    
    CONFIG2_DONE_q1 : SLE
      port map(D => CORECONFIGP_0_CONFIG2_DONE, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CONFIG2_DONE_q1\);
    
    CONFIG2_DONE_clk_base : SLE
      port map(D => \CONFIG2_DONE_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CONFIG2_DONE_clk_base\);
    
    CONFIG1_DONE_clk_base : SLE
      port map(D => \CONFIG1_DONE_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CONFIG1_DONE_clk_base\);
    
    sm0_areset_n_rcosc_RNIKFSA : CLKINT
      port map(A => sm0_areset_n_rcosc_0, Y => 
        \sm0_areset_n_rcosc\);
    
    mss_ready_select : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un6_fic_2_apb_m_preset_n_clk_base\, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_select\);
    
    un6_fic_2_apb_m_preset_n_clk_base : CFG2
      generic map(INIT => x"8")

      port map(A => \FIC_2_APB_M_PRESET_N_clk_base\, B => 
        \mss_ready_state\, Y => 
        \un6_fic_2_apb_m_preset_n_clk_base\);
    
    \count_ddr[4]\ : SLE
      port map(D => \count_ddr_s[4]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[4]_net_1\);
    
    \count_ddr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[6]_net_1\, S => \count_ddr_s[7]\, Y => 
        OPEN, FCO => \count_ddr_cry[7]_net_1\);
    
    release_sdif0_core : SLE
      port map(D => VCC_net_1, CLK => FABOSC_0_RCOSC_25_50MHZ_O2F, 
        EN => VCC_net_1, ALn => \sm0_areset_n_rcosc\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \release_sdif0_core\);
    
    POWER_ON_RESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => m2s010_som_sb_0_POWER_ON_RESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \POWER_ON_RESET_N_q1\);
    
    \count_ddr[12]\ : SLE
      port map(D => \count_ddr_s[12]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[12]_net_1\);
    
    ddr_settled : SLE
      port map(D => VCC_net_1, CLK => FABOSC_0_RCOSC_25_50MHZ_O2F, 
        EN => \un14_count_ddr\, ALn => \sm0_areset_n_rcosc\, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \ddr_settled\);
    
    \count_ddr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[8]_net_1\, S => \count_ddr_s[9]\, Y => 
        OPEN, FCO => \count_ddr_cry[9]_net_1\);
    
    \count_ddr[6]\ : SLE
      port map(D => \count_ddr_s[6]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[6]_net_1\);
    
    CONFIG1_DONE_q1 : SLE
      port map(D => CORECONFIGP_0_CONFIG1_DONE, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CONFIG1_DONE_q1\);
    
    un14_count_ddr_6 : CFG2
      generic map(INIT => x"1")

      port map(A => \count_ddr[6]_net_1\, B => 
        \count_ddr[7]_net_1\, Y => \un14_count_ddr_6\);
    
    sdif3_spll_lock_q1 : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => \sm0_areset_n_clk_base\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sdif3_spll_lock_q1\);
    
    release_sdif0_core_clk_base : SLE
      port map(D => \release_sdif0_core_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \release_sdif0_core_clk_base\);
    
    sdif3_spll_lock_q2 : SLE
      port map(D => \sdif3_spll_lock_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sdif3_spll_lock_q2\);
    
    RESET_N_M2F_clk_base : SLE
      port map(D => \RESET_N_M2F_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RESET_N_M2F_clk_base\);
    
    un1_next_ddr_ready_0_sqmuxa : CFG4
      generic map(INIT => x"F888")

      port map(A => \sdif3_spll_lock_q2\, B => 
        \sm0_state[3]_net_1\, C => \ddr_settled_clk_base\, D => 
        \sm0_state[2]_net_1\, Y => \un1_next_ddr_ready_0_sqmuxa\);
    
    \count_ddr[13]\ : SLE
      port map(D => \count_ddr_s[13]_net_1\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[13]_net_1\);
    
    \sm0_state_ns[5]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => \CONFIG2_DONE_clk_base\, B => 
        \sm0_state[1]_net_1\, C => \un8_ddr_settled_clk_base\, D
         => \sm0_state[2]_net_1\, Y => \sm0_state_ns[5]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_GPIO_6_IO is

    port( GPIO_6_PAD_0                      : inout std_logic := 'Z';
          GPIO_6_Y_0                        : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F_OE : in    std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F    : in    std_logic
        );

end m2s010_som_sb_GPIO_6_IO;

architecture DEF_ARCH of m2s010_som_sb_GPIO_6_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      generic map(IOSTD => "LVCMOS33")

      port map(PAD => GPIO_6_PAD_0, D => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F, E => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F_OE, Y => GPIO_6_Y_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreConfigP is

    port( CORECONFIGP_0_MDDR_APBmslave_PRDATA              : in    std_logic_vector(15 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR   : in    std_logic_vector(15 downto 2);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA  : out   std_logic_vector(17 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA  : in    std_logic_vector(16 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PWDATA              : out   std_logic_vector(15 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PADDR               : out   std_logic_vector(10 downto 2);
          CORECONFIGP_0_MDDR_APBmslave_PSLVERR             : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PSELx               : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx   : in    std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PREADY              : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PENABLE             : out   std_logic;
          INIT_DONE                                        : in    std_logic;
          CORECONFIGP_0_APB_S_PCLK_i                       : in    std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE  : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PWRITE              : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY  : out   std_logic;
          CORECONFIGP_0_CONFIG2_DONE                       : out   std_logic;
          CORECONFIGP_0_CONFIG1_DONE                       : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK                         : in    std_logic;
          CORECONFIGP_0_APB_S_PRESET_N                     : in    std_logic
        );

end CoreConfigP;

architecture DEF_ARCH of CoreConfigP is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \state_d[2]\, GND_net_1, \paddr[12]_net_1\, 
        \paddr_26\, \paddr[13]_net_1\, \paddr_27\, 
        \paddr[15]_net_1\, \paddr_29\, \soft_reset_reg[11]_net_1\, 
        \un17_int_psel\, \soft_reset_reg[12]_net_1\, 
        \soft_reset_reg[13]_net_1\, \soft_reset_reg[14]_net_1\, 
        \soft_reset_reg[15]_net_1\, \soft_reset_reg[16]_net_1\, 
        \CORECONFIGP_0_CONFIG1_DONE\, \un8_int_psel\, 
        \CORECONFIGP_0_CONFIG2_DONE\, \prdata[15]\, 
        \state[1]_net_1\, \prdata[16]\, \int_prdata_5_sqmuxa\, 
        \soft_reset_reg[0]_net_1\, \soft_reset_reg[1]_net_1\, 
        \soft_reset_reg[2]_net_1\, \soft_reset_reg[3]_net_1\, 
        \soft_reset_reg[4]_net_1\, \soft_reset_reg[5]_net_1\, 
        \soft_reset_reg[6]_net_1\, \soft_reset_reg[7]_net_1\, 
        \soft_reset_reg[8]_net_1\, \soft_reset_reg[9]_net_1\, 
        \soft_reset_reg[10]_net_1\, prdata_N_12_i, \prdata[1]\, 
        \prdata[2]\, \prdata[3]\, \prdata[4]\, \prdata[5]\, 
        \prdata[6]\, \prdata[7]\, \prdata[8]\, \prdata[9]\, 
        \prdata[10]\, \prdata[11]\, \prdata[12]\, \prdata[13]\, 
        \prdata[14]\, \FIC_2_APB_M_PREADY_0_RNO\, pslverr, 
        \state[0]_net_1\, \state_ns[0]\, \state_ns[1]\, \psel\, 
        \state_d_i[2]\, \INIT_DONE_q1\, \INIT_DONE_q2\, 
        \MDDR_PENABLE_0_1\, \soft_reset_reg_m_0[15]\, 
        \soft_reset_reg_m_0[3]\, \soft_reset_reg_m_0[11]\, 
        \soft_reset_reg_m_0[4]\, \soft_reset_reg_m_0[8]\, 
        \soft_reset_reg_m_0[13]\, \soft_reset_reg_m_0[12]\, 
        \soft_reset_reg_m_0[2]\, \soft_reset_reg_m_0[7]\, 
        \soft_reset_reg_m_0[14]\, \un20_int_psel\, 
        \soft_reset_reg_m_1[1]\, \soft_reset_reg_m[1]\, 
        un1_N_3_mux_0, \prdata_0_iv_1[16]_net_1\, 
        \int_prdata_4_sqmuxa\, \MDDR_PSEL_0_x\, pready, 
        un1_fic_2_apb_m_psel_i_0, \prdata_m11_0_a3_1\, 
        \prdata_m4_e\, INIT_DONE_q2_m_2_0, un6_m1_e_1, 
        \un11_int_psel\, \CORECONFIGP_0_MDDR_APBmslave_PSELx\, 
        prdata_m11_0_a3_0, \int_prdata_0_sqmuxa_a0\, 
        \prdata_0_iv_0_tz[5]_net_1\, \control_reg_1_m[1]\
         : std_logic;

begin 

    CORECONFIGP_0_MDDR_APBmslave_PSELx <= 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\;
    CORECONFIGP_0_CONFIG2_DONE <= \CORECONFIGP_0_CONFIG2_DONE\;
    CORECONFIGP_0_CONFIG1_DONE <= \CORECONFIGP_0_CONFIG1_DONE\;

    \soft_reset_reg[13]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(13), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[13]_net_1\);
    
    \pwdata[15]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(15), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(15));
    
    prdata_m11_0_a3_0_1 : CFG4
      generic map(INIT => x"135F")

      port map(A => \soft_reset_reg[0]_net_1\, B => 
        \CORECONFIGP_0_CONFIG1_DONE\, C => \un20_int_psel\, D => 
        \un11_int_psel\, Y => prdata_m11_0_a3_0);
    
    \pwdata[8]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(8), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(8));
    
    \prdata_0_iv_RNO[13]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), D => 
        \soft_reset_reg[13]_net_1\, Y => \soft_reset_reg_m_0[13]\);
    
    \pwdata[3]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(3), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(3));
    
    \soft_reset_reg[10]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(10), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[10]_net_1\);
    
    \prdata_0_iv[12]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => un1_N_3_mux_0, B => \soft_reset_reg_m_0[12]\, 
        C => CORECONFIGP_0_MDDR_APBmslave_PRDATA(12), D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[12]\);
    
    \paddr[8]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(8), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(8));
    
    \prdata_0_iv_RNO[14]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), D => 
        \soft_reset_reg[14]_net_1\, Y => \soft_reset_reg_m_0[14]\);
    
    \soft_reset_reg[2]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(2), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[2]_net_1\);
    
    \pwdata[5]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(5), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(5));
    
    \prdata_0_iv_RNO[2]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), D => 
        \soft_reset_reg[2]_net_1\, Y => \soft_reset_reg_m_0[2]\);
    
    \paddr[5]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(5), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(5));
    
    INIT_DONE_q1 : SLE
      port map(D => INIT_DONE, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => VCC_net_1, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \INIT_DONE_q1\);
    
    \FIC_2_APB_M_PRDATA_0[7]\ : SLE
      port map(D => \prdata[7]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(7));
    
    \paddr[3]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(3));
    
    \pwdata[9]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(9), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(9));
    
    \control_reg_1[0]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un8_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CORECONFIGP_0_CONFIG1_DONE\);
    
    \prdata_0_iv_1[16]\ : CFG3
      generic map(INIT => x"20")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), Y => 
        \prdata_0_iv_1[16]_net_1\);
    
    MDDR_PENABLE_0_1 : CFG4
      generic map(INIT => x"0100")

      port map(A => \paddr[12]_net_1\, B => \paddr[13]_net_1\, C
         => \paddr[15]_net_1\, D => \state[1]_net_1\, Y => 
        \MDDR_PENABLE_0_1\);
    
    \pwdata[7]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(7), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(7));
    
    FIC_2_APB_M_PREADY_0 : SLE
      port map(D => \state[1]_net_1\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => 
        \FIC_2_APB_M_PREADY_0_RNO\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY);
    
    \soft_reset_reg[9]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(9), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[9]_net_1\);
    
    \prdata_0_iv[16]\ : CFG4
      generic map(INIT => x"3320")

      port map(A => \soft_reset_reg[16]_net_1\, B => 
        un1_N_3_mux_0, C => \un20_int_psel\, D => 
        \prdata_0_iv_1[16]_net_1\, Y => \prdata[16]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \pwdata[1]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(1));
    
    \pwdata[13]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(13), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(13));
    
    \prdata_0_iv[11]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => un1_N_3_mux_0, B => \soft_reset_reg_m_0[11]\, 
        C => CORECONFIGP_0_MDDR_APBmslave_PRDATA(11), D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[11]\);
    
    \prdata_0_iv[10]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => \soft_reset_reg[10]_net_1\, B => 
        \int_prdata_4_sqmuxa\, C => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, D => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(10), Y => 
        \prdata[10]\);
    
    psel : SLE
      port map(D => \state_d_i[2]\, CLK => 
        CORECONFIGP_0_APB_S_PCLK_i, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => \psel\);
    
    \FIC_2_APB_M_PRDATA_0[17]\ : SLE
      port map(D => \int_prdata_5_sqmuxa\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(17));
    
    \FIC_2_APB_M_PRDATA_0[14]\ : SLE
      port map(D => \prdata[14]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(14));
    
    pwrite : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE);
    
    \pwdata[6]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(6), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(6));
    
    \paddr[12]\ : SLE
      port map(D => \paddr_26\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => VCC_net_1, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \paddr[12]_net_1\);
    
    int_prdata_5_sqmuxa : CFG4
      generic map(INIT => x"0020")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        un1_N_3_mux_0, C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), Y => 
        \int_prdata_5_sqmuxa\);
    
    \paddr[13]\ : SLE
      port map(D => \paddr_27\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => VCC_net_1, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \paddr[13]_net_1\);
    
    \FIC_2_APB_M_PRDATA_0[1]\ : SLE
      port map(D => \prdata[1]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(1));
    
    \prdata_0_iv_RNO_1[1]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \paddr[15]_net_1\, B => \paddr[13]_net_1\, Y
         => \soft_reset_reg_m_1[1]\);
    
    \prdata_0_iv[14]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => un1_N_3_mux_0, B => \soft_reset_reg_m_0[14]\, 
        C => CORECONFIGP_0_MDDR_APBmslave_PRDATA(14), D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[14]\);
    
    \soft_reset_reg[0]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[0]_net_1\);
    
    \pwdata[2]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(2), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(2));
    
    \prdata_0_iv[2]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => un1_N_3_mux_0, B => \soft_reset_reg_m_0[2]\, 
        C => CORECONFIGP_0_MDDR_APBmslave_PRDATA(2), D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[2]\);
    
    \state_ns_0[1]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \state[1]_net_1\, B => pready, C => 
        \state[0]_net_1\, Y => \state_ns[1]\);
    
    \prdata_0_iv[3]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => un1_N_3_mux_0, B => \soft_reset_reg_m_0[3]\, 
        C => CORECONFIGP_0_MDDR_APBmslave_PRDATA(3), D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[3]\);
    
    \FIC_2_APB_M_PRDATA_0[9]\ : SLE
      port map(D => \prdata[9]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(9));
    
    \prdata_0_iv_RNO[8]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), D => 
        \soft_reset_reg[8]_net_1\, Y => \soft_reset_reg_m_0[8]\);
    
    \FIC_2_APB_M_PRDATA_0[13]\ : SLE
      port map(D => \prdata[13]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(13));
    
    \soft_reset_reg[15]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(15), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[15]_net_1\);
    
    \paddr_RNINQ3R[13]\ : CFG3
      generic map(INIT => x"80")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, C => 
        \paddr[13]_net_1\, Y => un6_m1_e_1);
    
    \paddr[7]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(7), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(7));
    
    \FIC_2_APB_M_PRDATA_0[11]\ : SLE
      port map(D => \prdata[11]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(11));
    
    \prdata_0_iv[9]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => \soft_reset_reg[9]_net_1\, B => 
        \int_prdata_4_sqmuxa\, C => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, D => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(9), Y => \prdata[9]\);
    
    \prdata_0_iv[5]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => un1_N_3_mux_0, B => 
        \prdata_0_iv_0_tz[5]_net_1\, C => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(5), D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[5]\);
    
    \prdata_0_iv_RNO[3]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), D => 
        \soft_reset_reg[3]_net_1\, Y => \soft_reset_reg_m_0[3]\);
    
    \prdata_0_iv[13]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => un1_N_3_mux_0, B => \soft_reset_reg_m_0[13]\, 
        C => CORECONFIGP_0_MDDR_APBmslave_PRDATA(13), D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[13]\);
    
    \paddr[6]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(6), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(6));
    
    MDDR_PSEL_0 : CFG4
      generic map(INIT => x"0100")

      port map(A => \paddr[12]_net_1\, B => \paddr[13]_net_1\, C
         => \paddr[15]_net_1\, D => \psel\, Y => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\);
    
    \control_reg_1[1]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un8_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CORECONFIGP_0_CONFIG2_DONE\);
    
    \pwdata[11]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(11), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(11));
    
    \prdata_0_iv[15]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => un1_N_3_mux_0, B => \soft_reset_reg_m_0[15]\, 
        C => CORECONFIGP_0_MDDR_APBmslave_PRDATA(15), D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[15]\);
    
    \FIC_2_APB_M_PRDATA_0[2]\ : SLE
      port map(D => \prdata[2]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(2));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \soft_reset_reg[3]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(3), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[3]_net_1\);
    
    \soft_reset_reg[12]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(12), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[12]_net_1\);
    
    prdata_m11_0_a3_1_RNO : CFG2
      generic map(INIT => x"1")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), Y => 
        INIT_DONE_q2_m_2_0);
    
    \FIC_2_APB_M_PRDATA_0_RNO[0]\ : CFG3
      generic map(INIT => x"B1")

      port map(A => un1_N_3_mux_0, B => \prdata_m11_0_a3_1\, C
         => \prdata_m4_e\, Y => prdata_N_12_i);
    
    \FIC_2_APB_M_PRDATA_0[8]\ : SLE
      port map(D => \prdata[8]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(8));
    
    \state[0]\ : SLE
      port map(D => \state_ns[0]\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \state[0]_net_1\);
    
    un8_int_psel : CFG4
      generic map(INIT => x"0080")

      port map(A => un6_m1_e_1, B => \psel\, C => \un11_int_psel\, 
        D => \paddr[15]_net_1\, Y => \un8_int_psel\);
    
    prdata_m11_0_a3_0_0 : CFG3
      generic map(INIT => x"D0")

      port map(A => \paddr[13]_net_1\, B => \paddr[15]_net_1\, C
         => \psel\, Y => un1_N_3_mux_0);
    
    \prdata_0_iv[4]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => un1_N_3_mux_0, B => \soft_reset_reg_m_0[4]\, 
        C => CORECONFIGP_0_MDDR_APBmslave_PRDATA(4), D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[4]\);
    
    \FIC_2_APB_M_PRDATA_0[10]\ : SLE
      port map(D => \prdata[10]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(10));
    
    \pwdata[14]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(14), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(14));
    
    \prdata_0_iv_RNO[1]\ : CFG4
      generic map(INIT => x"8088")

      port map(A => \un20_int_psel\, B => 
        \soft_reset_reg[1]_net_1\, C => \soft_reset_reg_m_1[1]\, 
        D => \psel\, Y => \soft_reset_reg_m[1]\);
    
    \FIC_2_APB_M_PRDATA_0[16]\ : SLE
      port map(D => \prdata[16]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(16));
    
    \soft_reset_reg[4]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(4), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[4]_net_1\);
    
    FIC_2_APB_M_PSLVERR_0 : SLE
      port map(D => pslverr, CLK => CORECONFIGP_0_APB_S_PCLK, EN
         => \state[1]_net_1\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR);
    
    prdata_m11_0_a3_1 : CFG4
      generic map(INIT => x"70F0")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        INIT_DONE_q2_m_2_0, C => prdata_m11_0_a3_0, D => 
        \INIT_DONE_q2\, Y => \prdata_m11_0_a3_1\);
    
    \prdata_0_iv_RNO[7]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), D => 
        \soft_reset_reg[7]_net_1\, Y => \soft_reset_reg_m_0[7]\);
    
    state_s0_0_a2 : CFG2
      generic map(INIT => x"1")

      port map(A => \state[1]_net_1\, B => \state[0]_net_1\, Y
         => \state_d[2]\);
    
    \prdata_0_iv_RNO[12]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), D => 
        \soft_reset_reg[12]_net_1\, Y => \soft_reset_reg_m_0[12]\);
    
    \prdata_0_iv[1]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => \soft_reset_reg_m[1]\, B => 
        \control_reg_1_m[1]\, C => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, D => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(1), Y => \prdata[1]\);
    
    \soft_reset_reg[8]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(8), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[8]_net_1\);
    
    FIC_2_APB_M_PREADY_0_RNO : CFG4
      generic map(INIT => x"ECA0")

      port map(A => un1_fic_2_apb_m_psel_i_0, B => 
        \state[1]_net_1\, C => \state_d[2]\, D => pready, Y => 
        \FIC_2_APB_M_PREADY_0_RNO\);
    
    \prdata_0_iv[8]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => un1_N_3_mux_0, B => \soft_reset_reg_m_0[8]\, 
        C => CORECONFIGP_0_MDDR_APBmslave_PRDATA(8), D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[8]\);
    
    paddr_26 : CFG3
      generic map(INIT => x"D8")

      port map(A => \state_d[2]\, B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(12), C => 
        \paddr[12]_net_1\, Y => \paddr_26\);
    
    \FIC_2_APB_M_PRDATA_0[3]\ : SLE
      port map(D => \prdata[3]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(3));
    
    \prdata_0_iv_RNO[4]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), D => 
        \soft_reset_reg[4]_net_1\, Y => \soft_reset_reg_m_0[4]\);
    
    \prdata_0_iv[6]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => \soft_reset_reg[6]_net_1\, B => 
        \int_prdata_4_sqmuxa\, C => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, D => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(6), Y => \prdata[6]\);
    
    MDDR_PSEL_0_x_RNIH9T41 : CFG3
      generic map(INIT => x"DF")

      port map(A => \MDDR_PSEL_0_x\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PREADY, C => \psel\, Y => 
        pready);
    
    \pwdata[10]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(10), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(10));
    
    \prdata_0_iv[7]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => un1_N_3_mux_0, B => \soft_reset_reg_m_0[7]\, 
        C => CORECONFIGP_0_MDDR_APBmslave_PRDATA(7), D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[7]\);
    
    paddr_27 : CFG3
      generic map(INIT => x"D8")

      port map(A => \state_d[2]\, B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(13), C => 
        \paddr[13]_net_1\, Y => \paddr_27\);
    
    INIT_DONE_q2 : SLE
      port map(D => \INIT_DONE_q1\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INIT_DONE_q2\);
    
    \prdata_0_iv_0_tz[5]\ : CFG4
      generic map(INIT => x"0A40")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        \soft_reset_reg[5]_net_1\, C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), Y => 
        \prdata_0_iv_0_tz[5]_net_1\);
    
    \FIC_2_APB_M_PRDATA_0[0]\ : SLE
      port map(D => prdata_N_12_i, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(0));
    
    \state[1]\ : SLE
      port map(D => \state_ns[1]\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \state[1]_net_1\);
    
    \soft_reset_reg[6]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(6), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[6]_net_1\);
    
    \prdata_0_iv_RNO_0[1]\ : CFG4
      generic map(INIT => x"C0C8")

      port map(A => \un11_int_psel\, B => 
        \CORECONFIGP_0_CONFIG2_DONE\, C => 
        \int_prdata_0_sqmuxa_a0\, D => \psel\, Y => 
        \control_reg_1_m[1]\);
    
    FIC_2_APB_M_PSLVERR_0_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PSLVERR, B => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => pslverr);
    
    int_prdata_4_sqmuxa : CFG4
      generic map(INIT => x"7030")

      port map(A => \paddr[15]_net_1\, B => \psel\, C => 
        \un20_int_psel\, D => \paddr[13]_net_1\, Y => 
        \int_prdata_4_sqmuxa\);
    
    un20_int_psel : CFG3
      generic map(INIT => x"02")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), Y => 
        \un20_int_psel\);
    
    \soft_reset_reg[7]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(7), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[7]_net_1\);
    
    \soft_reset_reg[11]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(11), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[11]_net_1\);
    
    \paddr[4]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(4));
    
    int_prdata_0_sqmuxa_a0 : CFG3
      generic map(INIT => x"40")

      port map(A => \paddr[15]_net_1\, B => \un11_int_psel\, C
         => \paddr[13]_net_1\, Y => \int_prdata_0_sqmuxa_a0\);
    
    un11_int_psel : CFG3
      generic map(INIT => x"01")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), Y => 
        \un11_int_psel\);
    
    \pwdata[12]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(12), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(12));
    
    \paddr[9]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(9), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(9));
    
    \FIC_2_APB_M_PRDATA_0[15]\ : SLE
      port map(D => \prdata[15]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(15));
    
    un1_next_FIC_2_APB_M_PREADY_0_sqmuxa_0_a3 : CFG2
      generic map(INIT => x"8")

      port map(A => \state_d[2]\, B => un1_fic_2_apb_m_psel_i_0, 
        Y => \state_ns[0]\);
    
    \soft_reset_reg[1]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[1]_net_1\);
    
    prdata_m4_e : CFG4
      generic map(INIT => x"0100")

      port map(A => \paddr[12]_net_1\, B => \paddr[13]_net_1\, C
         => \paddr[15]_net_1\, D => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(0), Y => 
        \prdata_m4_e\);
    
    MDDR_PSEL_0_x : CFG3
      generic map(INIT => x"01")

      port map(A => \paddr[12]_net_1\, B => \paddr[13]_net_1\, C
         => \paddr[15]_net_1\, Y => \MDDR_PSEL_0_x\);
    
    \soft_reset_reg[16]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(16), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[16]_net_1\);
    
    \pwdata[0]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(0));
    
    \FIC_2_APB_M_PRDATA_0[4]\ : SLE
      port map(D => \prdata[4]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(4));
    
    \pwdata[4]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(4), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(4));
    
    MDDR_PENABLE_0 : SLE
      port map(D => \MDDR_PENABLE_0_1\, CLK => 
        CORECONFIGP_0_APB_S_PCLK_i, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE);
    
    \FIC_2_APB_M_PRDATA_0[12]\ : SLE
      port map(D => \prdata[12]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(12));
    
    \paddr[2]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(2));
    
    \paddr[10]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(10), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(10));
    
    state_s0_0_a2_i : CFG2
      generic map(INIT => x"E")

      port map(A => \state[1]_net_1\, B => \state[0]_net_1\, Y
         => \state_d_i[2]\);
    
    \prdata_0_iv_RNO[15]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), D => 
        \soft_reset_reg[15]_net_1\, Y => \soft_reset_reg_m_0[15]\);
    
    \FIC_2_APB_M_PRDATA_0[6]\ : SLE
      port map(D => \prdata[6]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(6));
    
    paddr_29 : CFG3
      generic map(INIT => x"D8")

      port map(A => \state_d[2]\, B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(15), C => 
        \paddr[15]_net_1\, Y => \paddr_29\);
    
    \soft_reset_reg[14]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(14), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[14]_net_1\);
    
    un17_int_psel : CFG4
      generic map(INIT => x"0080")

      port map(A => un6_m1_e_1, B => \psel\, C => \un20_int_psel\, 
        D => \paddr[15]_net_1\, Y => \un17_int_psel\);
    
    \prdata_0_iv_RNO[11]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), D => 
        \soft_reset_reg[11]_net_1\, Y => \soft_reset_reg_m_0[11]\);
    
    \paddr[15]\ : SLE
      port map(D => \paddr_29\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => VCC_net_1, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \paddr[15]_net_1\);
    
    un1_fic_2_apb_m_psel : CFG2
      generic map(INIT => x"4")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx, Y => 
        un1_fic_2_apb_m_psel_i_0);
    
    \soft_reset_reg[5]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(5), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[5]_net_1\);
    
    \FIC_2_APB_M_PRDATA_0[5]\ : SLE
      port map(D => \prdata[5]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(5));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_CCC_0_FCCC is

    port( m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : in    std_logic;
          FAB_CCC_LOCK                              : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz                 : out   std_logic
        );

end m2s010_som_sb_CCC_0_FCCC;

architecture DEF_ARCH of m2s010_som_sb_CCC_0_FCCC is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CCC

            generic (INIT:std_logic_vector(209 downto 0) := "00" & x"0000000000000000000000000000000000000000000000000000"; 
        VCOFREQUENCY:real := 0.0);

    port( Y0              : out   std_logic;
          Y1              : out   std_logic;
          Y2              : out   std_logic;
          Y3              : out   std_logic;
          PRDATA          : out   std_logic_vector(7 downto 0);
          LOCK            : out   std_logic;
          BUSY            : out   std_logic;
          CLK0            : in    std_logic := 'U';
          CLK1            : in    std_logic := 'U';
          CLK2            : in    std_logic := 'U';
          CLK3            : in    std_logic := 'U';
          NGMUX0_SEL      : in    std_logic := 'U';
          NGMUX1_SEL      : in    std_logic := 'U';
          NGMUX2_SEL      : in    std_logic := 'U';
          NGMUX3_SEL      : in    std_logic := 'U';
          NGMUX0_HOLD_N   : in    std_logic := 'U';
          NGMUX1_HOLD_N   : in    std_logic := 'U';
          NGMUX2_HOLD_N   : in    std_logic := 'U';
          NGMUX3_HOLD_N   : in    std_logic := 'U';
          NGMUX0_ARST_N   : in    std_logic := 'U';
          NGMUX1_ARST_N   : in    std_logic := 'U';
          NGMUX2_ARST_N   : in    std_logic := 'U';
          NGMUX3_ARST_N   : in    std_logic := 'U';
          PLL_BYPASS_N    : in    std_logic := 'U';
          PLL_ARST_N      : in    std_logic := 'U';
          PLL_POWERDOWN_N : in    std_logic := 'U';
          GPD0_ARST_N     : in    std_logic := 'U';
          GPD1_ARST_N     : in    std_logic := 'U';
          GPD2_ARST_N     : in    std_logic := 'U';
          GPD3_ARST_N     : in    std_logic := 'U';
          PRESET_N        : in    std_logic := 'U';
          PCLK            : in    std_logic := 'U';
          PSEL            : in    std_logic := 'U';
          PENABLE         : in    std_logic := 'U';
          PWRITE          : in    std_logic := 'U';
          PADDR           : in    std_logic_vector(7 downto 2) := (others => 'U');
          PWDATA          : in    std_logic_vector(7 downto 0) := (others => 'U');
          CLK0_PAD        : in    std_logic := 'U';
          CLK1_PAD        : in    std_logic := 'U';
          CLK2_PAD        : in    std_logic := 'U';
          CLK3_PAD        : in    std_logic := 'U';
          GL0             : out   std_logic;
          GL1             : out   std_logic;
          GL2             : out   std_logic;
          GL3             : out   std_logic;
          RCOSC_25_50MHZ  : in    std_logic := 'U';
          RCOSC_1MHZ      : in    std_logic := 'U';
          XTLOSC          : in    std_logic := 'U'
        );
  end component;

    signal GL0_net, VCC_net_1, GND_net_1 : std_logic;
    signal nc8, nc7, nc6, nc2, nc5, nc4, nc3, nc1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    GL0_INST : CLKINT
      port map(A => GL0_net, Y => m2s010_som_sb_0_CCC_71MHz);
    
    CCC_INST : CCC

              generic map(INIT => "00" & x"000007F88000044D64000318C6318C1F18C61E40404040404613",
         VCOFREQUENCY => 568.0)

      port map(Y0 => OPEN, Y1 => OPEN, Y2 => OPEN, Y3 => OPEN, 
        PRDATA(7) => nc8, PRDATA(6) => nc7, PRDATA(5) => nc6, 
        PRDATA(4) => nc2, PRDATA(3) => nc5, PRDATA(2) => nc4, 
        PRDATA(1) => nc3, PRDATA(0) => nc1, LOCK => FAB_CCC_LOCK, 
        BUSY => OPEN, CLK0 => VCC_net_1, CLK1 => VCC_net_1, CLK2
         => VCC_net_1, CLK3 => VCC_net_1, NGMUX0_SEL => GND_net_1, 
        NGMUX1_SEL => GND_net_1, NGMUX2_SEL => GND_net_1, 
        NGMUX3_SEL => GND_net_1, NGMUX0_HOLD_N => VCC_net_1, 
        NGMUX1_HOLD_N => VCC_net_1, NGMUX2_HOLD_N => VCC_net_1, 
        NGMUX3_HOLD_N => VCC_net_1, NGMUX0_ARST_N => VCC_net_1, 
        NGMUX1_ARST_N => VCC_net_1, NGMUX2_ARST_N => VCC_net_1, 
        NGMUX3_ARST_N => VCC_net_1, PLL_BYPASS_N => VCC_net_1, 
        PLL_ARST_N => VCC_net_1, PLL_POWERDOWN_N => VCC_net_1, 
        GPD0_ARST_N => VCC_net_1, GPD1_ARST_N => VCC_net_1, 
        GPD2_ARST_N => VCC_net_1, GPD3_ARST_N => VCC_net_1, 
        PRESET_N => GND_net_1, PCLK => VCC_net_1, PSEL => 
        VCC_net_1, PENABLE => VCC_net_1, PWRITE => VCC_net_1, 
        PADDR(7) => VCC_net_1, PADDR(6) => VCC_net_1, PADDR(5)
         => VCC_net_1, PADDR(4) => VCC_net_1, PADDR(3) => 
        VCC_net_1, PADDR(2) => VCC_net_1, PWDATA(7) => VCC_net_1, 
        PWDATA(6) => VCC_net_1, PWDATA(5) => VCC_net_1, PWDATA(4)
         => VCC_net_1, PWDATA(3) => VCC_net_1, PWDATA(2) => 
        VCC_net_1, PWDATA(1) => VCC_net_1, PWDATA(0) => VCC_net_1, 
        CLK0_PAD => GND_net_1, CLK1_PAD => GND_net_1, CLK2_PAD
         => GND_net_1, CLK3_PAD => GND_net_1, GL0 => GL0_net, GL1
         => OPEN, GL2 => OPEN, GL3 => OPEN, RCOSC_25_50MHZ => 
        GND_net_1, RCOSC_1MHZ => GND_net_1, XTLOSC => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_OTH_SPI_1_SS0_IO is

    port( SPI_1_SS0_OTH_0                      : inout std_logic := 'Z';
          OTH_SPI_1_SS0_Y_0                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F    : in    std_logic
        );

end m2s010_som_sb_OTH_SPI_1_SS0_IO;

architecture DEF_ARCH of m2s010_som_sb_OTH_SPI_1_SS0_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      port map(PAD => SPI_1_SS0_OTH_0, D => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F, E => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, Y => 
        OTH_SPI_1_SS0_Y_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_FABOSC_0_OSC is

    port( XTL                                       : in    std_logic;
          m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_O2F               : out   std_logic
        );

end m2s010_som_sb_FABOSC_0_OSC;

architecture DEF_ARCH of m2s010_som_sb_FABOSC_0_OSC is 

  component RCOSC_25_50MHZ_FAB
    port( A      : in    std_logic := 'U';
          CLKOUT : out   std_logic
        );
  end component;

  component RCOSC_25_50MHZ
    generic (FREQUENCY:real := 50.0);

    port( CLKOUT : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component XTLOSC
    generic (MODE:std_logic_vector(1 downto 0) := "11"; 
        FREQUENCY:real := 20.0);

    port( XTL    : in    std_logic := 'U';
          CLKOUT : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_RCOSC_25_50MHZ_CLKINT, N_RCOSC_25_50MHZ_CLKOUT, 
        GND_net_1, VCC_net_1 : std_logic;

begin 


    I_RCOSC_25_50MHZ_FAB : RCOSC_25_50MHZ_FAB
      port map(A => N_RCOSC_25_50MHZ_CLKOUT, CLKOUT => 
        N_RCOSC_25_50MHZ_CLKINT);
    
    I_RCOSC_25_50MHZ : RCOSC_25_50MHZ
      generic map(FREQUENCY => 50.0)

      port map(CLKOUT => N_RCOSC_25_50MHZ_CLKOUT);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    I_XTLOSC : XTLOSC
      generic map(MODE => "11", FREQUENCY => 20.0)

      port map(XTL => XTL, CLKOUT => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC);
    
    I_RCOSC_25_50MHZ_FAB_CLKINT : CLKINT
      port map(A => N_RCOSC_25_50MHZ_CLKINT, Y => 
        FABOSC_0_RCOSC_25_50MHZ_O2F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb is

    port( MDDR_DQS                                  : inout std_logic_vector(1 downto 0) := (others => 'Z');
          MDDR_DQ                                   : inout std_logic_vector(15 downto 0) := (others => 'Z');
          MDDR_DM_RDQS                              : inout std_logic_vector(1 downto 0) := (others => 'Z');
          MDDR_BA                                   : out   std_logic_vector(2 downto 0);
          MDDR_ADDR                                 : out   std_logic_vector(15 downto 0);
          CoreAPB3_0_APBmslave0_PADDR               : out   std_logic_vector(7 downto 0);
          m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR    : out   std_logic_vector(15 downto 12);
          CoreAPB3_0_APBmslave0_PWDATA              : out   std_logic_vector(7 downto 0);
          MAC_MII_TXD_c                             : out   std_logic_vector(3 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA_m            : in    std_logic_vector(7 downto 0);
          Y_net_0                                   : in    std_logic_vector(3 downto 0);
          MAC_MII_RXD_c                             : in    std_logic_vector(3 downto 0);
          SPI_1_SS0_OTH_0                           : inout std_logic := 'Z';
          DEBOUNCE_OUT_net_0_0                      : in    std_logic;
          GPIO_7_PADI_0                             : inout std_logic := 'Z';
          GPIO_6_PAD_0                              : inout std_logic := 'Z';
          GPIO_1_BI_0                               : inout std_logic := 'Z';
          SPI_1_SS0_CAM_0                           : inout std_logic := 'Z';
          SPI_1_CLK_0                               : inout std_logic := 'Z';
          SPI_0_SS1                                 : out   std_logic;
          SPI_0_SS0                                 : inout std_logic := 'Z';
          SPI_0_DO                                  : out   std_logic;
          SPI_0_DI                                  : in    std_logic;
          SPI_0_CLK                                 : inout std_logic := 'Z';
          MMUART_1_TXD                              : out   std_logic;
          MMUART_1_RXD                              : in    std_logic;
          MDDR_WE_N                                 : out   std_logic;
          MDDR_RESET_N                              : out   std_logic;
          MDDR_RAS_N                                : out   std_logic;
          MDDR_ODT                                  : out   std_logic;
          MDDR_DQS_TMATCH_0_OUT                     : out   std_logic;
          MDDR_DQS_TMATCH_0_IN                      : in    std_logic;
          MDDR_CS_N                                 : out   std_logic;
          MDDR_CKE                                  : out   std_logic;
          MDDR_CAS_N                                : out   std_logic;
          I2C_1_SDA                                 : inout std_logic := 'Z';
          I2C_1_SCL                                 : inout std_logic := 'Z';
          GPIO_31_BI                                : inout std_logic := 'Z';
          GPIO_26_BI                                : inout std_logic := 'Z';
          GPIO_25_BI                                : inout std_logic := 'Z';
          GPIO_20_OUT                               : out   std_logic;
          GPIO_18_BI                                : inout std_logic := 'Z';
          GPIO_17_BI                                : inout std_logic := 'Z';
          GPIO_16_BI                                : inout std_logic := 'Z';
          GPIO_15_BI                                : inout std_logic := 'Z';
          GPIO_14_BI                                : inout std_logic := 'Z';
          GPIO_12_BI                                : inout std_logic := 'Z';
          GPIO_4_BI                                 : inout std_logic := 'Z';
          GPIO_3_BI                                 : inout std_logic := 'Z';
          GPIO_0_BI                                 : inout std_logic := 'Z';
          CoreAPB3_0_APBmslave0_PENABLE             : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx    : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE              : out   std_logic;
          MAC_MII_MDC_c                             : out   std_logic;
          GPIO_22_M2F_c                             : out   std_logic;
          GPIO_21_M2F_c                             : out   std_logic;
          m2s010_som_sb_0_GPIO_28_SW_RESET          : out   std_logic;
          MMUART_0_TXD_M2F_c                        : out   std_logic;
          GPIO_24_M2F_c                             : out   std_logic;
          GPIO_5_M2F_c                              : out   std_logic;
          GPIO_8_M2F_c                              : out   std_logic;
          GPIO_11_M2F_c                             : out   std_logic;
          MAC_MII_TX_EN_c                           : out   std_logic;
          MAC_MII_COL_c                             : in    std_logic;
          MAC_MII_CRS_c                             : in    std_logic;
          CommsFPGA_top_0_INT                       : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY_i_m_i        : in    std_logic;
          DEBOUNCE_OUT_1_c                          : in    std_logic;
          DEBOUNCE_OUT_2_c                          : in    std_logic;
          MMUART_0_RXD_F2M_c                        : in    std_logic;
          MAC_MII_RX_CLK_c                          : in    std_logic;
          MAC_MII_RX_DV_c                           : in    std_logic;
          MAC_MII_RX_ER_c                           : in    std_logic;
          MAC_MII_TX_CLK_c                          : in    std_logic;
          MDDR_CLK_N                                : out   std_logic;
          MDDR_CLK                                  : out   std_logic;
          XTL                                       : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz                 : out   std_logic;
          m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : inout std_logic := 'Z';
          SPI_1_DI_CAM_c                            : in    std_logic;
          SPI_1_DI_OTH_c                            : in    std_logic;
          CommsFPGA_top_0_CAMERA_NODE               : in    std_logic;
          DEVRST_N                                  : in    std_logic;
          m2s010_som_sb_0_POWER_ON_RESET_N          : out   std_logic;
          MAC_MII_MDIO                              : inout std_logic := 'Z';
          SPI_1_DO_CAM_c                            : inout std_logic := 'Z';
          SPI_1_DO_OTH                              : out   std_logic
        );

end m2s010_som_sb;

architecture DEF_ARCH of m2s010_som_sb is 

  component m2s010_som_sb_GPIO_1_IO
    port( GPIO_1_BI_0                       : inout   std_logic;
          GPIO_1_in_0                       : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_1_M2F_OE : in    std_logic := 'U';
          GPIO_1_M2F                        : in    std_logic := 'U'
        );
  end component;

  component m2s010_som_sb_CAM_SPI_1_CLK_IO
    port( CAM_SPI_1_CLK_Y_0                    : out   std_logic;
          SPI_1_CLK_0                          : inout   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic := 'U';
          m2s010_som_sb_MSS_0_SPI_1_CLK_M2F    : in    std_logic := 'U'
        );
  end component;

  component m2s010_som_sb_GPIO_7_IO
    port( GPIO_7_PADI_0                     : inout   std_logic;
          GPIO_7_Y_0                        : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F_OE : in    std_logic := 'U';
          m2s010_som_sb_MSS_0_GPIO_7_M2F    : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component m2s010_som_sb_CAM_SPI_1_SS0_IO
    port( SPI_1_SS0_CAM_0                      : inout   std_logic;
          CAM_SPI_1_SS0_Y_0                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic := 'U';
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F    : in    std_logic := 'U'
        );
  end component;

  component m2s010_som_sb_MSS
    port( CORECONFIGP_0_MDDR_APBmslave_PWDATA              : in    std_logic_vector(15 downto 0) := (others => 'U');
          CORECONFIGP_0_MDDR_APBmslave_PADDR               : in    std_logic_vector(10 downto 2) := (others => 'U');
          MAC_MII_RXD_c                                    : in    std_logic_vector(3 downto 0) := (others => 'U');
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA  : in    std_logic_vector(17 downto 0) := (others => 'U');
          Y_net_0                                          : in    std_logic_vector(3 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PRDATA_m                   : in    std_logic_vector(7 downto 0) := (others => 'U');
          CORECONFIGP_0_MDDR_APBmslave_PRDATA              : out   std_logic_vector(15 downto 0);
          MAC_MII_TXD_c                                    : out   std_logic_vector(3 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA  : out   std_logic_vector(16 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR   : out   std_logic_vector(15 downto 2);
          CoreAPB3_0_APBmslave0_PWDATA                     : out   std_logic_vector(7 downto 0);
          m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR           : out   std_logic_vector(15 downto 12);
          CoreAPB3_0_APBmslave0_PADDR                      : out   std_logic_vector(7 downto 0);
          MDDR_ADDR                                        : out   std_logic_vector(15 downto 0);
          MDDR_BA                                          : out   std_logic_vector(2 downto 0);
          MDDR_DM_RDQS                                     : inout   std_logic_vector(1 downto 0);
          MDDR_DQ                                          : inout   std_logic_vector(15 downto 0);
          MDDR_DQS                                         : inout   std_logic_vector(1 downto 0);
          CAM_SPI_1_CLK_Y_0                                : in    std_logic := 'U';
          GPIO_7_Y_0                                       : in    std_logic := 'U';
          GPIO_6_Y_0                                       : in    std_logic := 'U';
          DEBOUNCE_OUT_net_0_0                             : in    std_logic := 'U';
          GPIO_1_in_0                                      : in    std_logic := 'U';
          MDDR_CLK                                         : out   std_logic;
          MDDR_CLK_N                                       : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PWRITE              : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PSELx               : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PENABLE             : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz                        : in    std_logic := 'U';
          MAC_MII_TX_CLK_c                                 : in    std_logic := 'U';
          SPI_1_SS0_MX_Y                                   : in    std_logic := 'U';
          SPI_1_DI                                         : in    std_logic := 'U';
          MAC_MII_RX_ER_c                                  : in    std_logic := 'U';
          MAC_MII_RX_DV_c                                  : in    std_logic := 'U';
          MAC_MII_RX_CLK_c                                 : in    std_logic := 'U';
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR : in    std_logic := 'U';
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY  : in    std_logic := 'U';
          MMUART_0_RXD_F2M_c                               : in    std_logic := 'U';
          DEBOUNCE_OUT_2_c                                 : in    std_logic := 'U';
          DEBOUNCE_OUT_1_c                                 : in    std_logic := 'U';
          BIBUF_0_Y                                        : in    std_logic := 'U';
          FAB_CCC_LOCK                                     : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY_i_m_i               : in    std_logic := 'U';
          CommsFPGA_top_0_INT                              : in    std_logic := 'U';
          MAC_MII_CRS_c                                    : in    std_logic := 'U';
          MAC_MII_COL_c                                    : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PSLVERR             : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PREADY              : out   std_logic;
          MAC_MII_TX_EN_c                                  : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE             : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F                : out   std_logic;
          SPI_1_DO_CAM_c                                   : out   std_logic;
          GPIO_11_M2F_c                                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_CLK_M2F                : out   std_logic;
          GPIO_8_M2F_c                                     : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F                   : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F_OE                : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F                   : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F_OE                : out   std_logic;
          GPIO_5_M2F_c                                     : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE  : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx   : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE : out   std_logic;
          GPIO_24_M2F_c                                    : out   std_logic;
          MMUART_0_TXD_M2F_c                               : out   std_logic;
          m2s010_som_sb_0_GPIO_28_SW_RESET                 : out   std_logic;
          GPIO_21_M2F_c                                    : out   std_logic;
          GPIO_22_M2F_c                                    : out   std_logic;
          m2s010_som_sb_MSS_0_MAC_MII_MDO                  : out   std_logic;
          m2s010_som_sb_MSS_0_MAC_MII_MDO_EN               : out   std_logic;
          MAC_MII_MDC_c                                    : out   std_logic;
          GPIO_1_M2F                                       : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_1_M2F_OE                : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F          : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE                     : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx           : out   std_logic;
          CoreAPB3_0_APBmslave0_PENABLE                    : out   std_logic;
          GPIO_0_BI                                        : inout   std_logic;
          GPIO_3_BI                                        : inout   std_logic;
          GPIO_4_BI                                        : inout   std_logic;
          GPIO_12_BI                                       : inout   std_logic;
          GPIO_14_BI                                       : inout   std_logic;
          GPIO_15_BI                                       : inout   std_logic;
          GPIO_16_BI                                       : inout   std_logic;
          GPIO_17_BI                                       : inout   std_logic;
          GPIO_18_BI                                       : inout   std_logic;
          GPIO_20_OUT                                      : out   std_logic;
          GPIO_25_BI                                       : inout   std_logic;
          GPIO_26_BI                                       : inout   std_logic;
          GPIO_31_BI                                       : inout   std_logic;
          I2C_1_SCL                                        : inout   std_logic;
          I2C_1_SDA                                        : inout   std_logic;
          MDDR_CAS_N                                       : out   std_logic;
          MDDR_CKE                                         : out   std_logic;
          MDDR_CS_N                                        : out   std_logic;
          MDDR_DQS_TMATCH_0_IN                             : in    std_logic := 'U';
          MDDR_DQS_TMATCH_0_OUT                            : out   std_logic;
          MDDR_ODT                                         : out   std_logic;
          MDDR_RAS_N                                       : out   std_logic;
          MDDR_RESET_N                                     : out   std_logic;
          MDDR_WE_N                                        : out   std_logic;
          MMUART_1_RXD                                     : in    std_logic := 'U';
          MMUART_1_TXD                                     : out   std_logic;
          SPI_0_CLK                                        : inout   std_logic;
          SPI_0_DI                                         : in    std_logic := 'U';
          SPI_0_DO                                         : out   std_logic;
          SPI_0_SS0                                        : inout   std_logic;
          SPI_0_SS1                                        : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK_i                       : out   std_logic;
          CORECONFIGP_0_APB_S_PRESET_N                     : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK                         : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CoreResetP
    port( CORECONFIGP_0_CONFIG2_DONE              : in    std_logic := 'U';
          CORECONFIGP_0_CONFIG1_DONE              : in    std_logic := 'U';
          CORECONFIGP_0_APB_S_PRESET_N            : in    std_logic := 'U';
          m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F : in    std_logic := 'U';
          m2s010_som_sb_0_POWER_ON_RESET_N        : in    std_logic := 'U';
          INIT_DONE                               : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_O2F             : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz               : in    std_logic := 'U'
        );
  end component;

  component SYSRESET
    port( POWER_ON_RESET_N : out   std_logic;
          DEVRST_N         : in    std_logic := 'U'
        );
  end component;

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component m2s010_som_sb_GPIO_6_IO
    port( GPIO_6_PAD_0                      : inout   std_logic;
          GPIO_6_Y_0                        : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F_OE : in    std_logic := 'U';
          m2s010_som_sb_MSS_0_GPIO_6_M2F    : in    std_logic := 'U'
        );
  end component;

  component CoreConfigP
    port( CORECONFIGP_0_MDDR_APBmslave_PRDATA              : in    std_logic_vector(15 downto 0) := (others => 'U');
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR   : in    std_logic_vector(15 downto 2) := (others => 'U');
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA  : out   std_logic_vector(17 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA  : in    std_logic_vector(16 downto 0) := (others => 'U');
          CORECONFIGP_0_MDDR_APBmslave_PWDATA              : out   std_logic_vector(15 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PADDR               : out   std_logic_vector(10 downto 2);
          CORECONFIGP_0_MDDR_APBmslave_PSLVERR             : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PSELx               : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx   : in    std_logic := 'U';
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PREADY              : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PENABLE             : out   std_logic;
          INIT_DONE                                        : in    std_logic := 'U';
          CORECONFIGP_0_APB_S_PCLK_i                       : in    std_logic := 'U';
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE  : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PWRITE              : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY  : out   std_logic;
          CORECONFIGP_0_CONFIG2_DONE                       : out   std_logic;
          CORECONFIGP_0_CONFIG1_DONE                       : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK                         : in    std_logic := 'U';
          CORECONFIGP_0_APB_S_PRESET_N                     : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component m2s010_som_sb_CCC_0_FCCC
    port( m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : in    std_logic := 'U';
          FAB_CCC_LOCK                              : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz                 : out   std_logic
        );
  end component;

  component m2s010_som_sb_OTH_SPI_1_SS0_IO
    port( SPI_1_SS0_OTH_0                      : inout   std_logic;
          OTH_SPI_1_SS0_Y_0                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic := 'U';
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F    : in    std_logic := 'U'
        );
  end component;

  component m2s010_som_sb_FABOSC_0_OSC
    port( XTL                                       : in    std_logic := 'U';
          m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_O2F               : out   std_logic
        );
  end component;

    signal BIBUF_0_Y, m2s010_som_sb_MSS_0_MAC_MII_MDO, 
        m2s010_som_sb_MSS_0_MAC_MII_MDO_EN, 
        \m2s010_som_sb_0_POWER_ON_RESET_N\, SPI_1_SS0_MX_Y, 
        \OTH_SPI_1_SS0_Y[0]\, \CAM_SPI_1_SS0_Y[0]\, SPI_1_DI, 
        \CAM_SPI_1_CLK_Y[0]\, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F, FAB_CCC_LOCK, 
        \m2s010_som_sb_0_CCC_71MHz\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[0]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[1]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[2]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[3]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[4]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[5]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[6]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[7]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[8]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[9]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[10]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[11]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[12]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[13]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[14]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[15]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[5]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[6]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[7]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[8]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[9]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[10]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[12]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[13]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[15]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[0]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[1]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[2]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[3]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[4]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[5]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[6]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[7]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[8]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[9]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[10]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[11]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[12]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[13]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[14]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[15]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[16]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[17]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[0]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[1]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[2]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[3]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[4]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[5]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[6]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[7]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[8]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[9]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[10]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[11]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[12]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[13]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[14]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[15]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[16]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[0]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[1]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[2]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[3]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[4]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[5]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[6]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[7]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[8]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[9]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[10]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[11]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[12]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[13]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[14]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[15]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[2]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[3]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[4]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[5]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[6]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[7]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[8]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[9]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR, 
        CORECONFIGP_0_MDDR_APBmslave_PSELx, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, 
        CORECONFIGP_0_MDDR_APBmslave_PREADY, 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE, INIT_DONE, 
        CORECONFIGP_0_APB_S_PCLK_i, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY, 
        CORECONFIGP_0_CONFIG2_DONE, CORECONFIGP_0_CONFIG1_DONE, 
        CORECONFIGP_0_APB_S_PCLK, CORECONFIGP_0_APB_S_PRESET_N, 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        FABOSC_0_RCOSC_25_50MHZ_O2F, \GPIO_1_in[0]\, 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE, GPIO_1_M2F, 
        \GPIO_6_Y[0]\, m2s010_som_sb_MSS_0_GPIO_6_M2F_OE, 
        m2s010_som_sb_MSS_0_GPIO_6_M2F, \GPIO_7_Y[0]\, 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE, 
        m2s010_som_sb_MSS_0_GPIO_7_M2F, GND_net_1, VCC_net_1
         : std_logic;
    signal nc2, nc4, nc3, nc1 : std_logic;

    for all : m2s010_som_sb_GPIO_1_IO
	Use entity work.m2s010_som_sb_GPIO_1_IO(DEF_ARCH);
    for all : m2s010_som_sb_CAM_SPI_1_CLK_IO
	Use entity work.m2s010_som_sb_CAM_SPI_1_CLK_IO(DEF_ARCH);
    for all : m2s010_som_sb_GPIO_7_IO
	Use entity work.m2s010_som_sb_GPIO_7_IO(DEF_ARCH);
    for all : m2s010_som_sb_CAM_SPI_1_SS0_IO
	Use entity work.m2s010_som_sb_CAM_SPI_1_SS0_IO(DEF_ARCH);
    for all : m2s010_som_sb_MSS
	Use entity work.m2s010_som_sb_MSS(DEF_ARCH);
    for all : CoreResetP
	Use entity work.CoreResetP(DEF_ARCH);
    for all : m2s010_som_sb_GPIO_6_IO
	Use entity work.m2s010_som_sb_GPIO_6_IO(DEF_ARCH);
    for all : CoreConfigP
	Use entity work.CoreConfigP(DEF_ARCH);
    for all : m2s010_som_sb_CCC_0_FCCC
	Use entity work.m2s010_som_sb_CCC_0_FCCC(DEF_ARCH);
    for all : m2s010_som_sb_OTH_SPI_1_SS0_IO
	Use entity work.m2s010_som_sb_OTH_SPI_1_SS0_IO(DEF_ARCH);
    for all : m2s010_som_sb_FABOSC_0_OSC
	Use entity work.m2s010_som_sb_FABOSC_0_OSC(DEF_ARCH);
begin 

    m2s010_som_sb_0_CCC_71MHz <= \m2s010_som_sb_0_CCC_71MHz\;
    m2s010_som_sb_0_POWER_ON_RESET_N <= 
        \m2s010_som_sb_0_POWER_ON_RESET_N\;

    GPIO_1 : m2s010_som_sb_GPIO_1_IO
      port map(GPIO_1_BI_0 => GPIO_1_BI_0, GPIO_1_in_0 => 
        \GPIO_1_in[0]\, m2s010_som_sb_MSS_0_GPIO_1_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE, GPIO_1_M2F => 
        GPIO_1_M2F);
    
    CAM_SPI_1_CLK : m2s010_som_sb_CAM_SPI_1_CLK_IO
      port map(CAM_SPI_1_CLK_Y_0 => \CAM_SPI_1_CLK_Y[0]\, 
        SPI_1_CLK_0 => SPI_1_CLK_0, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F => 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F);
    
    GPIO_7 : m2s010_som_sb_GPIO_7_IO
      port map(GPIO_7_PADI_0 => GPIO_7_PADI_0, GPIO_7_Y_0 => 
        \GPIO_7_Y[0]\, m2s010_som_sb_MSS_0_GPIO_7_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE, 
        m2s010_som_sb_MSS_0_GPIO_7_M2F => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    CAM_SPI_1_SS0 : m2s010_som_sb_CAM_SPI_1_SS0_IO
      port map(SPI_1_SS0_CAM_0 => SPI_1_SS0_CAM_0, 
        CAM_SPI_1_SS0_Y_0 => \CAM_SPI_1_SS0_Y[0]\, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F);
    
    m2s010_som_sb_MSS_0 : m2s010_som_sb_MSS
      port map(CORECONFIGP_0_MDDR_APBmslave_PWDATA(15) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(14) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[14]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(13) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[13]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(12) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[12]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(11) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[11]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(1) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[1]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(0) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[0]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[2]\, MAC_MII_RXD_c(3)
         => MAC_MII_RXD_c(3), MAC_MII_RXD_c(2) => 
        MAC_MII_RXD_c(2), MAC_MII_RXD_c(1) => MAC_MII_RXD_c(1), 
        MAC_MII_RXD_c(0) => MAC_MII_RXD_c(0), 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(17) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[17]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(16) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[16]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(14) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[14]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(11) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[11]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[2]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(1) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[1]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(0) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[0]\, 
        Y_net_0(3) => Y_net_0(3), Y_net_0(2) => Y_net_0(2), 
        Y_net_0(1) => Y_net_0(1), Y_net_0(0) => Y_net_0(0), 
        CoreAPB3_0_APBmslave0_PRDATA_m(7) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(7), 
        CoreAPB3_0_APBmslave0_PRDATA_m(6) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(6), 
        CoreAPB3_0_APBmslave0_PRDATA_m(5) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(5), 
        CoreAPB3_0_APBmslave0_PRDATA_m(4) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(4), 
        CoreAPB3_0_APBmslave0_PRDATA_m(3) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(3), 
        CoreAPB3_0_APBmslave0_PRDATA_m(2) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(2), 
        CoreAPB3_0_APBmslave0_PRDATA_m(1) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(1), 
        CoreAPB3_0_APBmslave0_PRDATA_m(0) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(0), 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(15) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(14) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[14]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(13) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[13]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(12) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[12]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(11) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[11]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(1) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[1]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(0) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[0]\, 
        MAC_MII_TXD_c(3) => MAC_MII_TXD_c(3), MAC_MII_TXD_c(2)
         => MAC_MII_TXD_c(2), MAC_MII_TXD_c(1) => 
        MAC_MII_TXD_c(1), MAC_MII_TXD_c(0) => MAC_MII_TXD_c(0), 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(16) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[16]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(14) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[14]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(11) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[11]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[2]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[1]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[0]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(14) => nc2, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(11) => nc4, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15), 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14), 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13), 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12), 
        CoreAPB3_0_APBmslave0_PADDR(7) => 
        CoreAPB3_0_APBmslave0_PADDR(7), 
        CoreAPB3_0_APBmslave0_PADDR(6) => 
        CoreAPB3_0_APBmslave0_PADDR(6), 
        CoreAPB3_0_APBmslave0_PADDR(5) => 
        CoreAPB3_0_APBmslave0_PADDR(5), 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        CoreAPB3_0_APBmslave0_PADDR(4), 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(3), 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        CoreAPB3_0_APBmslave0_PADDR(2), 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        CoreAPB3_0_APBmslave0_PADDR(1), 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        CoreAPB3_0_APBmslave0_PADDR(0), MDDR_ADDR(15) => 
        MDDR_ADDR(15), MDDR_ADDR(14) => MDDR_ADDR(14), 
        MDDR_ADDR(13) => MDDR_ADDR(13), MDDR_ADDR(12) => 
        MDDR_ADDR(12), MDDR_ADDR(11) => MDDR_ADDR(11), 
        MDDR_ADDR(10) => MDDR_ADDR(10), MDDR_ADDR(9) => 
        MDDR_ADDR(9), MDDR_ADDR(8) => MDDR_ADDR(8), MDDR_ADDR(7)
         => MDDR_ADDR(7), MDDR_ADDR(6) => MDDR_ADDR(6), 
        MDDR_ADDR(5) => MDDR_ADDR(5), MDDR_ADDR(4) => 
        MDDR_ADDR(4), MDDR_ADDR(3) => MDDR_ADDR(3), MDDR_ADDR(2)
         => MDDR_ADDR(2), MDDR_ADDR(1) => MDDR_ADDR(1), 
        MDDR_ADDR(0) => MDDR_ADDR(0), MDDR_BA(2) => MDDR_BA(2), 
        MDDR_BA(1) => MDDR_BA(1), MDDR_BA(0) => MDDR_BA(0), 
        MDDR_DM_RDQS(1) => MDDR_DM_RDQS(1), MDDR_DM_RDQS(0) => 
        MDDR_DM_RDQS(0), MDDR_DQ(15) => MDDR_DQ(15), MDDR_DQ(14)
         => MDDR_DQ(14), MDDR_DQ(13) => MDDR_DQ(13), MDDR_DQ(12)
         => MDDR_DQ(12), MDDR_DQ(11) => MDDR_DQ(11), MDDR_DQ(10)
         => MDDR_DQ(10), MDDR_DQ(9) => MDDR_DQ(9), MDDR_DQ(8) => 
        MDDR_DQ(8), MDDR_DQ(7) => MDDR_DQ(7), MDDR_DQ(6) => 
        MDDR_DQ(6), MDDR_DQ(5) => MDDR_DQ(5), MDDR_DQ(4) => 
        MDDR_DQ(4), MDDR_DQ(3) => MDDR_DQ(3), MDDR_DQ(2) => 
        MDDR_DQ(2), MDDR_DQ(1) => MDDR_DQ(1), MDDR_DQ(0) => 
        MDDR_DQ(0), MDDR_DQS(1) => MDDR_DQS(1), MDDR_DQS(0) => 
        MDDR_DQS(0), CAM_SPI_1_CLK_Y_0 => \CAM_SPI_1_CLK_Y[0]\, 
        GPIO_7_Y_0 => \GPIO_7_Y[0]\, GPIO_6_Y_0 => \GPIO_6_Y[0]\, 
        DEBOUNCE_OUT_net_0_0 => DEBOUNCE_OUT_net_0_0, GPIO_1_in_0
         => \GPIO_1_in[0]\, MDDR_CLK => MDDR_CLK, MDDR_CLK_N => 
        MDDR_CLK_N, CORECONFIGP_0_MDDR_APBmslave_PWRITE => 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE, 
        CORECONFIGP_0_MDDR_APBmslave_PSELx => 
        CORECONFIGP_0_MDDR_APBmslave_PSELx, 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE => 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE, 
        m2s010_som_sb_0_CCC_71MHz => \m2s010_som_sb_0_CCC_71MHz\, 
        MAC_MII_TX_CLK_c => MAC_MII_TX_CLK_c, SPI_1_SS0_MX_Y => 
        SPI_1_SS0_MX_Y, SPI_1_DI => SPI_1_DI, MAC_MII_RX_ER_c => 
        MAC_MII_RX_ER_c, MAC_MII_RX_DV_c => MAC_MII_RX_DV_c, 
        MAC_MII_RX_CLK_c => MAC_MII_RX_CLK_c, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY, 
        MMUART_0_RXD_F2M_c => MMUART_0_RXD_F2M_c, 
        DEBOUNCE_OUT_2_c => DEBOUNCE_OUT_2_c, DEBOUNCE_OUT_1_c
         => DEBOUNCE_OUT_1_c, BIBUF_0_Y => BIBUF_0_Y, 
        FAB_CCC_LOCK => FAB_CCC_LOCK, 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, CommsFPGA_top_0_INT
         => CommsFPGA_top_0_INT, MAC_MII_CRS_c => MAC_MII_CRS_c, 
        MAC_MII_COL_c => MAC_MII_COL_c, 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR => 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR, 
        CORECONFIGP_0_MDDR_APBmslave_PREADY => 
        CORECONFIGP_0_MDDR_APBmslave_PREADY, MAC_MII_TX_EN_c => 
        MAC_MII_TX_EN_c, m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F, SPI_1_DO_CAM_c => 
        SPI_1_DO_CAM_c, GPIO_11_M2F_c => GPIO_11_M2F_c, 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F => 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F, GPIO_8_M2F_c => 
        GPIO_8_M2F_c, m2s010_som_sb_MSS_0_GPIO_7_M2F => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F, 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE, 
        m2s010_som_sb_MSS_0_GPIO_6_M2F => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F, 
        m2s010_som_sb_MSS_0_GPIO_6_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F_OE, GPIO_5_M2F_c => 
        GPIO_5_M2F_c, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, 
        GPIO_24_M2F_c => GPIO_24_M2F_c, MMUART_0_TXD_M2F_c => 
        MMUART_0_TXD_M2F_c, m2s010_som_sb_0_GPIO_28_SW_RESET => 
        m2s010_som_sb_0_GPIO_28_SW_RESET, GPIO_21_M2F_c => 
        GPIO_21_M2F_c, GPIO_22_M2F_c => GPIO_22_M2F_c, 
        m2s010_som_sb_MSS_0_MAC_MII_MDO => 
        m2s010_som_sb_MSS_0_MAC_MII_MDO, 
        m2s010_som_sb_MSS_0_MAC_MII_MDO_EN => 
        m2s010_som_sb_MSS_0_MAC_MII_MDO_EN, MAC_MII_MDC_c => 
        MAC_MII_MDC_c, GPIO_1_M2F => GPIO_1_M2F, 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE, 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, GPIO_0_BI => GPIO_0_BI, 
        GPIO_3_BI => GPIO_3_BI, GPIO_4_BI => GPIO_4_BI, 
        GPIO_12_BI => GPIO_12_BI, GPIO_14_BI => GPIO_14_BI, 
        GPIO_15_BI => GPIO_15_BI, GPIO_16_BI => GPIO_16_BI, 
        GPIO_17_BI => GPIO_17_BI, GPIO_18_BI => GPIO_18_BI, 
        GPIO_20_OUT => GPIO_20_OUT, GPIO_25_BI => GPIO_25_BI, 
        GPIO_26_BI => GPIO_26_BI, GPIO_31_BI => GPIO_31_BI, 
        I2C_1_SCL => I2C_1_SCL, I2C_1_SDA => I2C_1_SDA, 
        MDDR_CAS_N => MDDR_CAS_N, MDDR_CKE => MDDR_CKE, MDDR_CS_N
         => MDDR_CS_N, MDDR_DQS_TMATCH_0_IN => 
        MDDR_DQS_TMATCH_0_IN, MDDR_DQS_TMATCH_0_OUT => 
        MDDR_DQS_TMATCH_0_OUT, MDDR_ODT => MDDR_ODT, MDDR_RAS_N
         => MDDR_RAS_N, MDDR_RESET_N => MDDR_RESET_N, MDDR_WE_N
         => MDDR_WE_N, MMUART_1_RXD => MMUART_1_RXD, MMUART_1_TXD
         => MMUART_1_TXD, SPI_0_CLK => SPI_0_CLK, SPI_0_DI => 
        SPI_0_DI, SPI_0_DO => SPI_0_DO, SPI_0_SS0 => SPI_0_SS0, 
        SPI_0_SS1 => SPI_0_SS1, CORECONFIGP_0_APB_S_PCLK_i => 
        CORECONFIGP_0_APB_S_PCLK_i, CORECONFIGP_0_APB_S_PRESET_N
         => CORECONFIGP_0_APB_S_PRESET_N, 
        CORECONFIGP_0_APB_S_PCLK => CORECONFIGP_0_APB_S_PCLK);
    
    SPI_1_SS0_MX : MX2
      port map(A => \OTH_SPI_1_SS0_Y[0]\, B => 
        \CAM_SPI_1_SS0_Y[0]\, S => CommsFPGA_top_0_CAMERA_NODE, Y
         => SPI_1_SS0_MX_Y);
    
    CORERESETP_0 : CoreResetP
      port map(CORECONFIGP_0_CONFIG2_DONE => 
        CORECONFIGP_0_CONFIG2_DONE, CORECONFIGP_0_CONFIG1_DONE
         => CORECONFIGP_0_CONFIG1_DONE, 
        CORECONFIGP_0_APB_S_PRESET_N => 
        CORECONFIGP_0_APB_S_PRESET_N, 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        m2s010_som_sb_0_POWER_ON_RESET_N => 
        \m2s010_som_sb_0_POWER_ON_RESET_N\, INIT_DONE => 
        INIT_DONE, FABOSC_0_RCOSC_25_50MHZ_O2F => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, m2s010_som_sb_0_CCC_71MHz
         => \m2s010_som_sb_0_CCC_71MHz\);
    
    SYSRESET_POR : SYSRESET
      port map(POWER_ON_RESET_N => 
        \m2s010_som_sb_0_POWER_ON_RESET_N\, DEVRST_N => DEVRST_N);
    
    BIBUF_0 : BIBUF
      port map(PAD => MAC_MII_MDIO, D => 
        m2s010_som_sb_MSS_0_MAC_MII_MDO, E => 
        m2s010_som_sb_MSS_0_MAC_MII_MDO_EN, Y => BIBUF_0_Y);
    
    SPI_1_D0_OUT : OUTBUF
      port map(D => SPI_1_DO_CAM_c, PAD => SPI_1_DO_OTH);
    
    GPIO_6 : m2s010_som_sb_GPIO_6_IO
      port map(GPIO_6_PAD_0 => GPIO_6_PAD_0, GPIO_6_Y_0 => 
        \GPIO_6_Y[0]\, m2s010_som_sb_MSS_0_GPIO_6_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F_OE, 
        m2s010_som_sb_MSS_0_GPIO_6_M2F => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F);
    
    CORECONFIGP_0 : CoreConfigP
      port map(CORECONFIGP_0_MDDR_APBmslave_PRDATA(15) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(14) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[14]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(13) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[13]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(12) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[12]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(11) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[11]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(1) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[1]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(0) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[0]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(14) => nc3, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(11) => nc1, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(17) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[17]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(16) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[16]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(14) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[14]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(11) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[11]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[2]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(1) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[1]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(0) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[0]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(16) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[16]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(14) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[14]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(11) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[11]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[2]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[1]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[0]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(15) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(14) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[14]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(13) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[13]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(12) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[12]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(11) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[11]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(1) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[1]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(0) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[0]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR => 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR, 
        CORECONFIGP_0_MDDR_APBmslave_PSELx => 
        CORECONFIGP_0_MDDR_APBmslave_PSELx, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, 
        CORECONFIGP_0_MDDR_APBmslave_PREADY => 
        CORECONFIGP_0_MDDR_APBmslave_PREADY, 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE => 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE, INIT_DONE => 
        INIT_DONE, CORECONFIGP_0_APB_S_PCLK_i => 
        CORECONFIGP_0_APB_S_PCLK_i, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE => 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY, 
        CORECONFIGP_0_CONFIG2_DONE => CORECONFIGP_0_CONFIG2_DONE, 
        CORECONFIGP_0_CONFIG1_DONE => CORECONFIGP_0_CONFIG1_DONE, 
        CORECONFIGP_0_APB_S_PCLK => CORECONFIGP_0_APB_S_PCLK, 
        CORECONFIGP_0_APB_S_PRESET_N => 
        CORECONFIGP_0_APB_S_PRESET_N);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    CCC_0 : m2s010_som_sb_CCC_0_FCCC
      port map(m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC, FAB_CCC_LOCK
         => FAB_CCC_LOCK, m2s010_som_sb_0_CCC_71MHz => 
        \m2s010_som_sb_0_CCC_71MHz\);
    
    SPI_1_DI_MX : MX2
      port map(A => SPI_1_DI_OTH_c, B => SPI_1_DI_CAM_c, S => 
        CommsFPGA_top_0_CAMERA_NODE, Y => SPI_1_DI);
    
    OTH_SPI_1_SS0 : m2s010_som_sb_OTH_SPI_1_SS0_IO
      port map(SPI_1_SS0_OTH_0 => SPI_1_SS0_OTH_0, 
        OTH_SPI_1_SS0_Y_0 => \OTH_SPI_1_SS0_Y[0]\, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F);
    
    FABOSC_0 : m2s010_som_sb_FABOSC_0_OSC
      port map(XTL => XTL, 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC, 
        FABOSC_0_RCOSC_25_50MHZ_O2F => 
        FABOSC_0_RCOSC_25_50MHZ_O2F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Debounce_1 is

    port( DEBOUNCE_IN_c_0  : in    std_logic;
          N_480            : in    std_logic;
          DEBOUNCE_OUT_2_c : out   std_logic;
          N_480_set        : in    std_logic;
          BIT_CLK          : in    std_logic
        );

end Debounce_1;

architecture DEF_ARCH of Debounce_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \debounce_cntr[1]_net_1\, VCC_net_1, 
        un2_debounce_in_i, un3_debounce_cntr_1_cry_1_S_1, 
        GND_net_1, \debounce_cntr[2]_net_1\, 
        un3_debounce_cntr_1_cry_2_S_1, \debounce_cntr[3]_net_1\, 
        un3_debounce_cntr_1_cry_3_S_1, \debounce_cntrrs[4]\, 
        un3_debounce_in_rs_1, \debounce_cntr[4]\, 
        un3_debounce_in_i, un3_debounce_cntr_1_cry_4_S_1, 
        \debounce_cntrrs[6]\, \debounce_cntr[6]\, 
        un3_debounce_cntr_1_cry_6_S_1, \debounce_cntr[5]\, 
        un3_debounce_cntr_1_cry_5_S_1, \debounce_cntr[7]\, 
        un3_debounce_cntr_1_cry_7_S_1, \debounce_cntrrs[8]\, 
        \debounce_cntr[8]_net_1\, un3_debounce_cntr_1_cry_8_S_1, 
        \debounce_cntrrs[9]\, \debounce_cntr[9]_net_1\, 
        un3_debounce_cntr_1_cry_9_S_1, \debounce_cntr[10]_net_1\, 
        un3_debounce_cntr_1_cry_10_S_1, \debounce_cntr[11]_net_1\, 
        un3_debounce_cntr_1_cry_11_S_1, \debounce_cntr[12]_net_1\, 
        un3_debounce_cntr_1_cry_12_S_1, \debounce_cntr[13]_net_1\, 
        un3_debounce_cntr_1_cry_13_S_1, \debounce_cntrrs[14]\, 
        \debounce_cntr[14]_net_1\, un3_debounce_cntr_1_cry_14_S_1, 
        \debounce_cntrrs[15]\, \debounce_cntr[15]_net_1\, 
        un3_debounce_cntr_1_s_15_S_1, \debounce_cntr[0]_net_1\, 
        \debounce_cntr_4[0]_net_1\, DEBOUNCE_OUT_2_crs, 
        un1_debounce_cntr, un3_debounce_cntr_1_s_1_274_FCO, 
        \un3_debounce_cntr_1_cry_1\, \un3_debounce_cntr_1_cry_2\, 
        \un3_debounce_cntr_1_cry_3\, \un3_debounce_cntr_1_cry_4\, 
        \un3_debounce_cntr_1_cry_5\, \un3_debounce_cntr_1_cry_6\, 
        \un3_debounce_cntr_1_cry_7\, \un3_debounce_cntr_1_cry_8\, 
        \un3_debounce_cntr_1_cry_9\, \un3_debounce_cntr_1_cry_10\, 
        \un3_debounce_cntr_1_cry_11\, 
        \un3_debounce_cntr_1_cry_12\, 
        \un3_debounce_cntr_1_cry_13\, 
        \un3_debounce_cntr_1_cry_14\, un1_debounce_cntr_11, 
        un1_debounce_cntr_10, un1_debounce_cntr_9, 
        un1_debounce_cntr_8 : std_logic;

begin 


    \debounce_cntr_0_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_5_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[5]\);
    
    un3_debounce_cntr_1_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[9]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_8\, S => 
        un3_debounce_cntr_1_cry_9_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_9\);
    
    \debounce_cntr_0_RNI48RR[0]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[4]\, B => 
        un3_debounce_in_rs_1, C => N_480_set, Y => 
        \debounce_cntr[4]\);
    
    \debounce_cntr[12]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_12_S_1, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un2_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[12]_net_1\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_8\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \debounce_cntr[9]_net_1\, B => 
        \debounce_cntr[8]_net_1\, C => \debounce_cntr[6]\, D => 
        \debounce_cntr[4]\, Y => un1_debounce_cntr_8);
    
    \DEBOUNCE_PROC.un3_debounce_in_rs\ : SLE
      port map(D => VCC_net_1, CLK => N_480, EN => VCC_net_1, ALn
         => un3_debounce_in_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => VCC_net_1, Q => 
        un3_debounce_in_rs_1);
    
    \debounce_cntr[15]\ : SLE
      port map(D => un3_debounce_cntr_1_s_15_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[15]\);
    
    un3_debounce_cntr_1_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_4\, S => 
        un3_debounce_cntr_1_cry_5_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_5\);
    
    un3_debounce_cntr_1_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[2]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_1\, S => 
        un3_debounce_cntr_1_cry_2_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_2\);
    
    \debounce_cntr[3]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_3_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[3]_net_1\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_9\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \debounce_cntr[2]_net_1\, B => 
        \debounce_cntr[1]_net_1\, C => \debounce_cntr[15]_net_1\, 
        D => \debounce_cntr[14]_net_1\, Y => un1_debounce_cntr_9);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_10\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[10]_net_1\, B => 
        \debounce_cntr[7]\, C => \debounce_cntr[5]\, D => 
        \debounce_cntr[3]_net_1\, Y => un1_debounce_cntr_10);
    
    debounce_out : SLE
      port map(D => un1_debounce_cntr, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un3_debounce_in_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => DEBOUNCE_OUT_2_crs);
    
    \debounce_cntr[10]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_10_S_1, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un2_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[10]_net_1\);
    
    un3_debounce_cntr_1_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_3\, S => 
        un3_debounce_cntr_1_cry_4_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_4\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \debounce_cntr[13]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_13_S_1, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un2_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[13]_net_1\);
    
    un3_debounce_cntr_1_cry_14 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[14]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_13\, S => 
        un3_debounce_cntr_1_cry_14_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_14\);
    
    \debounce_cntr_0_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_7_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[7]\);
    
    \debounce_cntr_RNIAJL01[14]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[14]\, B => 
        un3_debounce_in_rs_1, C => N_480_set, Y => 
        \debounce_cntr[14]_net_1\);
    
    un3_debounce_cntr_1_cry_13 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[13]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_12\, S => 
        un3_debounce_cntr_1_cry_13_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_13\);
    
    \debounce_cntr[9]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_9_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[9]\);
    
    un3_debounce_cntr_1_s_1_274 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[0]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un3_debounce_cntr_1_s_1_274_FCO);
    
    un3_debounce_cntr_1_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_6\, S => 
        un3_debounce_cntr_1_cry_7_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_7\);
    
    \debounce_cntr_RNIBKL01[15]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[15]\, B => 
        un3_debounce_in_rs_1, C => N_480_set, Y => 
        \debounce_cntr[15]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \DEBOUNCE_PROC.un2_debounce_in\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_480, B => DEBOUNCE_IN_c_0, Y => 
        un2_debounce_in_i);
    
    \debounce_cntr[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_1_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[1]_net_1\);
    
    \debounce_cntr_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_4_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[4]\);
    
    \debounce_cntr_RNIUINK[9]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[9]\, B => 
        un3_debounce_in_rs_1, C => N_480_set, Y => 
        \debounce_cntr[9]_net_1\);
    
    \debounce_cntr[14]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_14_S_1, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un3_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[14]\);
    
    un3_debounce_cntr_1_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_5\, S => 
        un3_debounce_cntr_1_cry_6_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_6\);
    
    un3_debounce_cntr_1_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[11]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_10\, S => 
        un3_debounce_cntr_1_cry_11_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_11\);
    
    \debounce_cntr_4[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => un1_debounce_cntr, B => 
        \debounce_cntr[0]_net_1\, Y => \debounce_cntr_4[0]_net_1\);
    
    \debounce_cntr[8]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_8_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[8]\);
    
    \debounce_cntr[0]\ : SLE
      port map(D => \debounce_cntr_4[0]_net_1\, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[0]_net_1\);
    
    \debounce_cntr_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_6_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[6]\);
    
    un3_debounce_cntr_1_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[8]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_7\, S => 
        un3_debounce_cntr_1_cry_8_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_8\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr\ : CFG4
      generic map(INIT => x"8000")

      port map(A => un1_debounce_cntr_11, B => 
        un1_debounce_cntr_10, C => un1_debounce_cntr_8, D => 
        un1_debounce_cntr_9, Y => un1_debounce_cntr);
    
    un3_debounce_cntr_1_cry_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[12]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_11\, S => 
        un3_debounce_cntr_1_cry_12_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_12\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_11\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[13]_net_1\, B => 
        \debounce_cntr[12]_net_1\, C => \debounce_cntr[11]_net_1\, 
        D => \debounce_cntr[0]_net_1\, Y => un1_debounce_cntr_11);
    
    un3_debounce_cntr_1_s_15 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[15]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_14\, S => 
        un3_debounce_cntr_1_s_15_S_1, Y => OPEN, FCO => OPEN);
    
    un3_debounce_cntr_1_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[10]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_9\, S => 
        un3_debounce_cntr_1_cry_10_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_10\);
    
    debounce_out_RNIEEKQ : CFG3
      generic map(INIT => x"F8")

      port map(A => un3_debounce_in_rs_1, B => N_480_set, C => 
        DEBOUNCE_OUT_2_crs, Y => DEBOUNCE_OUT_2_c);
    
    \debounce_cntr[2]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_2_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[2]_net_1\);
    
    \debounce_cntr[11]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_11_S_1, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un2_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[11]_net_1\);
    
    \debounce_cntr_0_RNI59RR[1]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[6]\, B => 
        un3_debounce_in_rs_1, C => N_480_set, Y => 
        \debounce_cntr[6]\);
    
    un3_debounce_cntr_1_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[1]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        un3_debounce_cntr_1_s_1_274_FCO, S => 
        un3_debounce_cntr_1_cry_1_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_1\);
    
    \debounce_cntr_RNITHNK[8]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[8]\, B => 
        un3_debounce_in_rs_1, C => N_480_set, Y => 
        \debounce_cntr[8]_net_1\);
    
    un3_debounce_cntr_1_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[3]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_2\, S => 
        un3_debounce_cntr_1_cry_3_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_3\);
    
    \DEBOUNCE_PROC.un3_debounce_in\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_480, B => DEBOUNCE_IN_c_0, Y => 
        un3_debounce_in_i);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Debounce_0 is

    port( DEBOUNCE_IN_c_0  : in    std_logic;
          N_480            : in    std_logic;
          DEBOUNCE_OUT_1_c : out   std_logic;
          N_480_set        : in    std_logic;
          BIT_CLK          : in    std_logic
        );

end Debounce_0;

architecture DEF_ARCH of Debounce_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \debounce_cntr[1]_net_1\, VCC_net_1, 
        un2_debounce_in_i, un3_debounce_cntr_1_cry_1_S_0, 
        GND_net_1, \debounce_cntr[2]_net_1\, 
        un3_debounce_cntr_1_cry_2_S_0, \debounce_cntr[3]_net_1\, 
        un3_debounce_cntr_1_cry_3_S_0, \debounce_cntrrs[4]\, 
        un3_debounce_in_rs_0, \debounce_cntr[4]\, 
        un3_debounce_in_i, un3_debounce_cntr_1_cry_4_S_0, 
        \debounce_cntrrs[6]\, \debounce_cntr[6]\, 
        un3_debounce_cntr_1_cry_6_S_0, \debounce_cntr[5]\, 
        un3_debounce_cntr_1_cry_5_S_0, \debounce_cntr[7]\, 
        un3_debounce_cntr_1_cry_7_S_0, \debounce_cntrrs[8]\, 
        \debounce_cntr[8]_net_1\, un3_debounce_cntr_1_cry_8_S_0, 
        \debounce_cntrrs[9]\, \debounce_cntr[9]_net_1\, 
        un3_debounce_cntr_1_cry_9_S_0, \debounce_cntr[10]_net_1\, 
        un3_debounce_cntr_1_cry_10_S_0, \debounce_cntr[11]_net_1\, 
        un3_debounce_cntr_1_cry_11_S_0, \debounce_cntr[12]_net_1\, 
        un3_debounce_cntr_1_cry_12_S_0, \debounce_cntr[13]_net_1\, 
        un3_debounce_cntr_1_cry_13_S_0, \debounce_cntrrs[14]\, 
        \debounce_cntr[14]_net_1\, un3_debounce_cntr_1_cry_14_S_0, 
        \debounce_cntrrs[15]\, \debounce_cntr[15]_net_1\, 
        un3_debounce_cntr_1_s_15_S_0, \debounce_cntr[0]_net_1\, 
        \debounce_cntr_4[0]_net_1\, DEBOUNCE_OUT_1_crs, 
        un1_debounce_cntr, un3_debounce_cntr_1_s_1_273_FCO, 
        \un3_debounce_cntr_1_cry_1\, \un3_debounce_cntr_1_cry_2\, 
        \un3_debounce_cntr_1_cry_3\, \un3_debounce_cntr_1_cry_4\, 
        \un3_debounce_cntr_1_cry_5\, \un3_debounce_cntr_1_cry_6\, 
        \un3_debounce_cntr_1_cry_7\, \un3_debounce_cntr_1_cry_8\, 
        \un3_debounce_cntr_1_cry_9\, \un3_debounce_cntr_1_cry_10\, 
        \un3_debounce_cntr_1_cry_11\, 
        \un3_debounce_cntr_1_cry_12\, 
        \un3_debounce_cntr_1_cry_13\, 
        \un3_debounce_cntr_1_cry_14\, un1_debounce_cntr_11, 
        un1_debounce_cntr_10, un1_debounce_cntr_9, 
        un1_debounce_cntr_8 : std_logic;

begin 


    \debounce_cntr_0_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_5_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[5]\);
    
    un3_debounce_cntr_1_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[9]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_8\, S => 
        un3_debounce_cntr_1_cry_9_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_9\);
    
    \debounce_cntr[12]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_12_S_0, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un2_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[12]_net_1\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_8\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \debounce_cntr[9]_net_1\, B => 
        \debounce_cntr[8]_net_1\, C => \debounce_cntr[6]\, D => 
        \debounce_cntr[4]\, Y => un1_debounce_cntr_8);
    
    \DEBOUNCE_PROC.un3_debounce_in_rs\ : SLE
      port map(D => VCC_net_1, CLK => N_480, EN => VCC_net_1, ALn
         => un3_debounce_in_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => VCC_net_1, Q => 
        un3_debounce_in_rs_0);
    
    \debounce_cntr_RNIRLFV[8]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => N_480_set, B => \debounce_cntrrs[8]\, C => 
        un3_debounce_in_rs_0, Y => \debounce_cntr[8]_net_1\);
    
    \debounce_cntr[15]\ : SLE
      port map(D => un3_debounce_cntr_1_s_15_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[15]\);
    
    un3_debounce_cntr_1_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_4\, S => 
        un3_debounce_cntr_1_cry_5_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_5\);
    
    un3_debounce_cntr_1_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[2]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_1\, S => 
        un3_debounce_cntr_1_cry_2_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_2\);
    
    \debounce_cntr[3]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_3_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[3]_net_1\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_9\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \debounce_cntr[2]_net_1\, B => 
        \debounce_cntr[1]_net_1\, C => \debounce_cntr[15]_net_1\, 
        D => \debounce_cntr[14]_net_1\, Y => un1_debounce_cntr_9);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_10\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[10]_net_1\, B => 
        \debounce_cntr[7]\, C => \debounce_cntr[5]\, D => 
        \debounce_cntr[3]_net_1\, Y => un1_debounce_cntr_10);
    
    debounce_out : SLE
      port map(D => un1_debounce_cntr, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un3_debounce_in_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => DEBOUNCE_OUT_1_crs);
    
    \debounce_cntr[10]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_10_S_0, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un2_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[10]_net_1\);
    
    un3_debounce_cntr_1_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_3\, S => 
        un3_debounce_cntr_1_cry_4_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_4\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \debounce_cntr[13]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_13_S_0, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un2_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[13]_net_1\);
    
    un3_debounce_cntr_1_cry_14 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[14]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_13\, S => 
        un3_debounce_cntr_1_cry_14_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_14\);
    
    \debounce_cntr_0_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_7_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[7]\);
    
    \debounce_cntr_RNI9NN31[15]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => N_480_set, B => \debounce_cntrrs[15]\, C => 
        un3_debounce_in_rs_0, Y => \debounce_cntr[15]_net_1\);
    
    un3_debounce_cntr_1_cry_13 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[13]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_12\, S => 
        un3_debounce_cntr_1_cry_13_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_13\);
    
    \debounce_cntr[9]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_9_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[9]\);
    
    un3_debounce_cntr_1_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_6\, S => 
        un3_debounce_cntr_1_cry_7_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_7\);
    
    \debounce_cntr_0_RNI3B611[1]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => N_480_set, B => \debounce_cntrrs[6]\, C => 
        un3_debounce_in_rs_0, Y => \debounce_cntr[6]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \DEBOUNCE_PROC.un2_debounce_in\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_480, B => DEBOUNCE_IN_c_0, Y => 
        un2_debounce_in_i);
    
    \debounce_cntr[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_1_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[1]_net_1\);
    
    \debounce_cntr_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_4_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[4]\);
    
    \debounce_cntr_RNI8MN31[14]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => N_480_set, B => \debounce_cntrrs[14]\, C => 
        un3_debounce_in_rs_0, Y => \debounce_cntr[14]_net_1\);
    
    \debounce_cntr[14]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_14_S_0, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un3_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[14]\);
    
    un3_debounce_cntr_1_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_5\, S => 
        un3_debounce_cntr_1_cry_6_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_6\);
    
    un3_debounce_cntr_1_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[11]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_10\, S => 
        un3_debounce_cntr_1_cry_11_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_11\);
    
    \debounce_cntr_RNISMFV[9]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => N_480_set, B => \debounce_cntrrs[9]\, C => 
        un3_debounce_in_rs_0, Y => \debounce_cntr[9]_net_1\);
    
    \debounce_cntr_4[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => un1_debounce_cntr, B => 
        \debounce_cntr[0]_net_1\, Y => \debounce_cntr_4[0]_net_1\);
    
    \debounce_cntr[8]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_8_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[8]\);
    
    \debounce_cntr[0]\ : SLE
      port map(D => \debounce_cntr_4[0]_net_1\, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[0]_net_1\);
    
    \debounce_cntr_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_6_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[6]\);
    
    un3_debounce_cntr_1_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[8]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_7\, S => 
        un3_debounce_cntr_1_cry_8_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_8\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr\ : CFG4
      generic map(INIT => x"8000")

      port map(A => un1_debounce_cntr_11, B => 
        un1_debounce_cntr_10, C => un1_debounce_cntr_8, D => 
        un1_debounce_cntr_9, Y => un1_debounce_cntr);
    
    un3_debounce_cntr_1_cry_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[12]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_11\, S => 
        un3_debounce_cntr_1_cry_12_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_12\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_11\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[13]_net_1\, B => 
        \debounce_cntr[12]_net_1\, C => \debounce_cntr[11]_net_1\, 
        D => \debounce_cntr[0]_net_1\, Y => un1_debounce_cntr_11);
    
    \debounce_cntr_0_RNI2A611[0]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => N_480_set, B => \debounce_cntrrs[4]\, C => 
        un3_debounce_in_rs_0, Y => \debounce_cntr[4]\);
    
    un3_debounce_cntr_1_s_15 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[15]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_14\, S => 
        un3_debounce_cntr_1_s_15_S_0, Y => OPEN, FCO => OPEN);
    
    un3_debounce_cntr_1_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[10]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_9\, S => 
        un3_debounce_cntr_1_cry_10_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_10\);
    
    \debounce_cntr[2]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_2_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[2]_net_1\);
    
    \debounce_cntr[11]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_11_S_0, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un2_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[11]_net_1\);
    
    un3_debounce_cntr_1_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[1]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        un3_debounce_cntr_1_s_1_273_FCO, S => 
        un3_debounce_cntr_1_cry_1_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_1\);
    
    debounce_out_RNICMQR : CFG3
      generic map(INIT => x"EA")

      port map(A => DEBOUNCE_OUT_1_crs, B => un3_debounce_in_rs_0, 
        C => N_480_set, Y => DEBOUNCE_OUT_1_c);
    
    un3_debounce_cntr_1_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[3]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_2\, S => 
        un3_debounce_cntr_1_cry_3_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_3\);
    
    un3_debounce_cntr_1_s_1_273 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[0]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un3_debounce_cntr_1_s_1_273_FCO);
    
    \DEBOUNCE_PROC.un3_debounce_in\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_480, B => DEBOUNCE_IN_c_0, Y => 
        un3_debounce_in_i);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Debounce is

    port( DEBOUNCE_IN_c_0      : in    std_logic;
          DEBOUNCE_OUT_net_0_0 : out   std_logic;
          N_480                : in    std_logic;
          N_480_set            : in    std_logic;
          BIT_CLK              : in    std_logic
        );

end Debounce;

architecture DEF_ARCH of Debounce is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \debounce_cntr[1]_net_1\, VCC_net_1, 
        un2_debounce_in_i, un3_debounce_cntr_1_cry_1_S, GND_net_1, 
        \debounce_cntr[2]_net_1\, un3_debounce_cntr_1_cry_2_S, 
        \debounce_cntr[3]_net_1\, un3_debounce_cntr_1_cry_3_S, 
        \debounce_cntrrs[4]\, un3_debounce_in_rs, 
        \debounce_cntr[4]\, un3_debounce_in_i, 
        un3_debounce_cntr_1_cry_4_S, \debounce_cntrrs[6]\, 
        \debounce_cntr[6]\, un3_debounce_cntr_1_cry_6_S, 
        \debounce_cntr[5]\, un3_debounce_cntr_1_cry_5_S, 
        \debounce_cntr[7]\, un3_debounce_cntr_1_cry_7_S, 
        \debounce_cntrrs[8]\, \debounce_cntr[8]_net_1\, 
        un3_debounce_cntr_1_cry_8_S, \debounce_cntrrs[9]\, 
        \debounce_cntr[9]_net_1\, un3_debounce_cntr_1_cry_9_S, 
        \debounce_cntr[10]_net_1\, un3_debounce_cntr_1_cry_10_S, 
        \debounce_cntr[11]_net_1\, un3_debounce_cntr_1_cry_11_S, 
        \debounce_cntr[12]_net_1\, un3_debounce_cntr_1_cry_12_S, 
        \debounce_cntr[13]_net_1\, un3_debounce_cntr_1_cry_13_S, 
        \debounce_cntrrs[14]\, \debounce_cntr[14]_net_1\, 
        un3_debounce_cntr_1_cry_14_S, \debounce_cntrrs[15]\, 
        \debounce_cntr[15]_net_1\, un3_debounce_cntr_1_s_15_S, 
        \debounce_cntr[0]_net_1\, \debounce_cntr_4[0]_net_1\, 
        \DEBOUNCE_OUT_net_0rs[0]\, un1_debounce_cntr, 
        un3_debounce_cntr_1_s_1_272_FCO, 
        \un3_debounce_cntr_1_cry_1\, \un3_debounce_cntr_1_cry_2\, 
        \un3_debounce_cntr_1_cry_3\, \un3_debounce_cntr_1_cry_4\, 
        \un3_debounce_cntr_1_cry_5\, \un3_debounce_cntr_1_cry_6\, 
        \un3_debounce_cntr_1_cry_7\, \un3_debounce_cntr_1_cry_8\, 
        \un3_debounce_cntr_1_cry_9\, \un3_debounce_cntr_1_cry_10\, 
        \un3_debounce_cntr_1_cry_11\, 
        \un3_debounce_cntr_1_cry_12\, 
        \un3_debounce_cntr_1_cry_13\, 
        \un3_debounce_cntr_1_cry_14\, un1_debounce_cntr_11, 
        un1_debounce_cntr_10, un1_debounce_cntr_9, 
        un1_debounce_cntr_8 : std_logic;

begin 


    \debounce_cntr_0_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_5_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[5]\);
    
    un3_debounce_cntr_1_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[9]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_8\, S => 
        un3_debounce_cntr_1_cry_9_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_9\);
    
    \debounce_cntr[12]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_12_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[12]_net_1\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_8\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \debounce_cntr[9]_net_1\, B => 
        \debounce_cntr[8]_net_1\, C => \debounce_cntr[6]\, D => 
        \debounce_cntr[4]\, Y => un1_debounce_cntr_8);
    
    \DEBOUNCE_PROC.un3_debounce_in_rs\ : SLE
      port map(D => VCC_net_1, CLK => N_480, EN => VCC_net_1, ALn
         => un3_debounce_in_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => VCC_net_1, Q => 
        un3_debounce_in_rs);
    
    \debounce_cntr[15]\ : SLE
      port map(D => un3_debounce_cntr_1_s_15_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[15]\);
    
    un3_debounce_cntr_1_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_4\, S => 
        un3_debounce_cntr_1_cry_5_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_5\);
    
    un3_debounce_cntr_1_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[2]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_1\, S => 
        un3_debounce_cntr_1_cry_2_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_2\);
    
    \debounce_cntr[3]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_3_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[3]_net_1\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_9\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \debounce_cntr[2]_net_1\, B => 
        \debounce_cntr[1]_net_1\, C => \debounce_cntr[15]_net_1\, 
        D => \debounce_cntr[14]_net_1\, Y => un1_debounce_cntr_9);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_10\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[10]_net_1\, B => 
        \debounce_cntr[7]\, C => \debounce_cntr[5]\, D => 
        \debounce_cntr[3]_net_1\, Y => un1_debounce_cntr_10);
    
    debounce_out : SLE
      port map(D => un1_debounce_cntr, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un3_debounce_in_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \DEBOUNCE_OUT_net_0rs[0]\);
    
    \debounce_cntr[10]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_10_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[10]_net_1\);
    
    un3_debounce_cntr_1_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_3\, S => 
        un3_debounce_cntr_1_cry_4_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_4\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \debounce_cntr_0_RNI0CHM[0]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => N_480_set, B => \debounce_cntrrs[4]\, C => 
        un3_debounce_in_rs, Y => \debounce_cntr[4]\);
    
    \debounce_cntr[13]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_13_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[13]_net_1\);
    
    un3_debounce_cntr_1_cry_14 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[14]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_13\, S => 
        un3_debounce_cntr_1_cry_14_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_14\);
    
    \debounce_cntr_0_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_7_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[7]\);
    
    \debounce_cntr_RNIPP7Q[8]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => N_480_set, B => \debounce_cntrrs[8]\, C => 
        un3_debounce_in_rs, Y => \debounce_cntr[8]_net_1\);
    
    un3_debounce_cntr_1_cry_13 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[13]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_12\, S => 
        un3_debounce_cntr_1_cry_13_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_13\);
    
    \debounce_cntr[9]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_9_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[9]\);
    
    \debounce_cntr_RNIQQ7Q[9]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => N_480_set, B => \debounce_cntrrs[9]\, C => 
        un3_debounce_in_rs, Y => \debounce_cntr[9]_net_1\);
    
    un3_debounce_cntr_1_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_6\, S => 
        un3_debounce_cntr_1_cry_7_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_7\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \DEBOUNCE_PROC.un2_debounce_in\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_480, B => DEBOUNCE_IN_c_0, Y => 
        un2_debounce_in_i);
    
    \debounce_cntr[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_1_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[1]_net_1\);
    
    \debounce_cntr_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_4_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[4]\);
    
    \debounce_cntr[14]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_14_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[14]\);
    
    un3_debounce_cntr_1_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_5\, S => 
        un3_debounce_cntr_1_cry_6_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_6\);
    
    un3_debounce_cntr_1_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[11]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_10\, S => 
        un3_debounce_cntr_1_cry_11_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_11\);
    
    \debounce_cntr_4[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => un1_debounce_cntr, B => 
        \debounce_cntr[0]_net_1\, Y => \debounce_cntr_4[0]_net_1\);
    
    \debounce_cntr_RNI7QPM[15]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => N_480_set, B => \debounce_cntrrs[15]\, C => 
        un3_debounce_in_rs, Y => \debounce_cntr[15]_net_1\);
    
    \debounce_cntr[8]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_8_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[8]\);
    
    \debounce_cntr[0]\ : SLE
      port map(D => \debounce_cntr_4[0]_net_1\, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[0]_net_1\);
    
    \debounce_cntr_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_6_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[6]\);
    
    debounce_out_RNIAU0T : CFG3
      generic map(INIT => x"EA")

      port map(A => \DEBOUNCE_OUT_net_0rs[0]\, B => 
        un3_debounce_in_rs, C => N_480_set, Y => 
        DEBOUNCE_OUT_net_0_0);
    
    un3_debounce_cntr_1_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[8]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_7\, S => 
        un3_debounce_cntr_1_cry_8_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_8\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr\ : CFG4
      generic map(INIT => x"8000")

      port map(A => un1_debounce_cntr_11, B => 
        un1_debounce_cntr_10, C => un1_debounce_cntr_8, D => 
        un1_debounce_cntr_9, Y => un1_debounce_cntr);
    
    un3_debounce_cntr_1_cry_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[12]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_11\, S => 
        un3_debounce_cntr_1_cry_12_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_12\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_11\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[13]_net_1\, B => 
        \debounce_cntr[12]_net_1\, C => \debounce_cntr[11]_net_1\, 
        D => \debounce_cntr[0]_net_1\, Y => un1_debounce_cntr_11);
    
    un3_debounce_cntr_1_s_15 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[15]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_14\, S => 
        un3_debounce_cntr_1_s_15_S, Y => OPEN, FCO => OPEN);
    
    un3_debounce_cntr_1_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[10]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_9\, S => 
        un3_debounce_cntr_1_cry_10_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_10\);
    
    un3_debounce_cntr_1_s_1_272 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[0]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un3_debounce_cntr_1_s_1_272_FCO);
    
    \debounce_cntr_RNI6PPM[14]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => N_480_set, B => \debounce_cntrrs[14]\, C => 
        un3_debounce_in_rs, Y => \debounce_cntr[14]_net_1\);
    
    \debounce_cntr[2]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_2_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[2]_net_1\);
    
    \debounce_cntr[11]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_11_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[11]_net_1\);
    
    \debounce_cntr_0_RNI1DHM[1]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => N_480_set, B => \debounce_cntrrs[6]\, C => 
        un3_debounce_in_rs, Y => \debounce_cntr[6]\);
    
    un3_debounce_cntr_1_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[1]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        un3_debounce_cntr_1_s_1_272_FCO, S => 
        un3_debounce_cntr_1_cry_1_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_1\);
    
    un3_debounce_cntr_1_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[3]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_2\, S => 
        un3_debounce_cntr_1_cry_3_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_3\);
    
    \DEBOUNCE_PROC.un3_debounce_in\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_480, B => DEBOUNCE_IN_c_0, Y => 
        un3_debounce_in_i);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity TriDebounce is

    port( DEBOUNCE_IN_c        : in    std_logic_vector(2 downto 0);
          DEBOUNCE_OUT_net_0_0 : out   std_logic;
          DEBOUNCE_OUT_2_c     : out   std_logic;
          DEBOUNCE_OUT_1_c     : out   std_logic;
          BIT_CLK              : in    std_logic;
          N_480_set            : in    std_logic;
          N_480                : in    std_logic
        );

end TriDebounce;

architecture DEF_ARCH of TriDebounce is 

  component Debounce_1
    port( DEBOUNCE_IN_c_0  : in    std_logic := 'U';
          N_480            : in    std_logic := 'U';
          DEBOUNCE_OUT_2_c : out   std_logic;
          N_480_set        : in    std_logic := 'U';
          BIT_CLK          : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component Debounce_0
    port( DEBOUNCE_IN_c_0  : in    std_logic := 'U';
          N_480            : in    std_logic := 'U';
          DEBOUNCE_OUT_1_c : out   std_logic;
          N_480_set        : in    std_logic := 'U';
          BIT_CLK          : in    std_logic := 'U'
        );
  end component;

  component Debounce
    port( DEBOUNCE_IN_c_0      : in    std_logic := 'U';
          DEBOUNCE_OUT_net_0_0 : out   std_logic;
          N_480                : in    std_logic := 'U';
          N_480_set            : in    std_logic := 'U';
          BIT_CLK              : in    std_logic := 'U'
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : Debounce_1
	Use entity work.Debounce_1(DEF_ARCH);
    for all : Debounce_0
	Use entity work.Debounce_0(DEF_ARCH);
    for all : Debounce
	Use entity work.Debounce(DEF_ARCH);
begin 


    DEBOUNCE_2_INST : Debounce_1
      port map(DEBOUNCE_IN_c_0 => DEBOUNCE_IN_c(2), N_480 => 
        N_480, DEBOUNCE_OUT_2_c => DEBOUNCE_OUT_2_c, N_480_set
         => N_480_set, BIT_CLK => BIT_CLK);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    DEBOUNCE_1_INST : Debounce_0
      port map(DEBOUNCE_IN_c_0 => DEBOUNCE_IN_c(1), N_480 => 
        N_480, DEBOUNCE_OUT_1_c => DEBOUNCE_OUT_1_c, N_480_set
         => N_480_set, BIT_CLK => BIT_CLK);
    
    DEBOUNCE_0_INST : Debounce
      port map(DEBOUNCE_IN_c_0 => DEBOUNCE_IN_c(0), 
        DEBOUNCE_OUT_net_0_0 => DEBOUNCE_OUT_net_0_0, N_480 => 
        N_480, N_480_set => N_480_set, BIT_CLK => BIT_CLK);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CRC16_Generator_0 is

    port( tx_crc_data : out   std_logic_vector(15 downto 0);
          N_518       : in    std_logic;
          N_519       : in    std_logic;
          N_228       : in    std_logic;
          N_520       : in    std_logic;
          N_521       : in    std_logic;
          N_516       : in    std_logic;
          N_517       : in    std_logic;
          N_522       : in    std_logic;
          tx_crc_gen  : in    std_logic;
          byte_clk_en : in    std_logic;
          BIT_CLK     : in    std_logic;
          N_9_0_i_i   : in    std_logic
        );

end CRC16_Generator_0;

architecture DEF_ARCH of CRC16_Generator_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \tx_crc_data[13]\, GND_net_1, \tx_crc_data[5]\, 
        \lfsr_q_0_sqmuxa\, VCC_net_1, \tx_crc_data[14]\, 
        \tx_crc_data[6]\, \tx_crc_data[15]\, \lfsr_c[15]\, 
        \tx_crc_data[0]\, \lfsr_c[0]\, \tx_crc_data[1]\, 
        \lfsr_c[1]\, \tx_crc_data[2]\, N_192_i, \tx_crc_data[3]\, 
        N_200_i, \tx_crc_data[4]\, N_195_i, N_201_i, N_193_i, 
        \tx_crc_data[7]\, N_194_i, \tx_crc_data[8]\, N_202_i_i, 
        \tx_crc_data[9]\, \lfsr_c[9]\, \tx_crc_data[10]\, 
        \tx_crc_data[11]\, \tx_crc_data[12]\, N_161_i
         : std_logic;

begin 

    tx_crc_data(15) <= \tx_crc_data[15]\;
    tx_crc_data(14) <= \tx_crc_data[14]\;
    tx_crc_data(13) <= \tx_crc_data[13]\;
    tx_crc_data(12) <= \tx_crc_data[12]\;
    tx_crc_data(11) <= \tx_crc_data[11]\;
    tx_crc_data(10) <= \tx_crc_data[10]\;
    tx_crc_data(9) <= \tx_crc_data[9]\;
    tx_crc_data(8) <= \tx_crc_data[8]\;
    tx_crc_data(7) <= \tx_crc_data[7]\;
    tx_crc_data(6) <= \tx_crc_data[6]\;
    tx_crc_data(5) <= \tx_crc_data[5]\;
    tx_crc_data(4) <= \tx_crc_data[4]\;
    tx_crc_data(3) <= \tx_crc_data[3]\;
    tx_crc_data(2) <= \tx_crc_data[2]\;
    tx_crc_data(1) <= \tx_crc_data[1]\;
    tx_crc_data(0) <= \tx_crc_data[0]\;

    \lfsr_q[9]\ : SLE
      port map(D => \lfsr_c[9]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => N_9_0_i_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_crc_data[9]\);
    
    \lfsr_c_0_a2_2_x2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[9]\, B => \tx_crc_data[8]\, C
         => N_517, D => N_516, Y => N_192_i);
    
    \lfsr_q[6]\ : SLE
      port map(D => N_193_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => N_9_0_i_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_crc_data[6]\);
    
    \lfsr_q[3]\ : SLE
      port map(D => N_200_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => N_9_0_i_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_crc_data[3]\);
    
    \lfsr_c_0_a2_2_x2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[13]\, B => \tx_crc_data[12]\, C
         => N_521, D => N_520, Y => N_193_i);
    
    \lfsr_q[10]\ : SLE
      port map(D => \tx_crc_data[2]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => N_9_0_i_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_crc_data[10]\);
    
    \lfsr_q[2]\ : SLE
      port map(D => N_192_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => N_9_0_i_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_crc_data[2]\);
    
    \lfsr_c_0_a2_0_x2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[14]\, B => \tx_crc_data[13]\, C
         => N_521, D => N_228, Y => N_194_i);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \lfsr_q[1]\ : SLE
      port map(D => \lfsr_c[1]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => N_9_0_i_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_crc_data[1]\);
    
    \lfsr_q[7]\ : SLE
      port map(D => N_194_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => N_9_0_i_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_crc_data[7]\);
    
    \lfsr_c_0_a2_0_x2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[10]\, B => \tx_crc_data[9]\, C
         => N_518, D => N_517, Y => N_200_i);
    
    \lfsr_q[4]\ : SLE
      port map(D => N_195_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => N_9_0_i_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_crc_data[4]\);
    
    \lfsr_q[11]\ : SLE
      port map(D => \tx_crc_data[3]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => N_9_0_i_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_crc_data[11]\);
    
    \lfsr_q[5]\ : SLE
      port map(D => N_201_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => N_9_0_i_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_crc_data[5]\);
    
    \lfsr_c_0_a2[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => N_161_i, B => \tx_crc_data[1]\, Y => 
        \lfsr_c[9]\);
    
    \lfsr_c_0_a2[1]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => N_194_i, B => N_200_i, C => N_161_i, D => 
        N_201_i, Y => \lfsr_c[1]\);
    
    \lfsr_q[0]\ : SLE
      port map(D => \lfsr_c[0]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => N_9_0_i_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_crc_data[0]\);
    
    \lfsr_c_0_a2[15]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => N_516, B => \lfsr_c[1]\, C => 
        \tx_crc_data[7]\, D => \tx_crc_data[8]\, Y => 
        \lfsr_c[15]\);
    
    \lfsr_q[12]\ : SLE
      port map(D => \tx_crc_data[4]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => N_9_0_i_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_crc_data[12]\);
    
    lfsr_q_0_sqmuxa : CFG2
      generic map(INIT => x"8")

      port map(A => byte_clk_en, B => tx_crc_gen, Y => 
        \lfsr_q_0_sqmuxa\);
    
    \lfsr_q[14]\ : SLE
      port map(D => \tx_crc_data[6]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => N_9_0_i_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_crc_data[14]\);
    
    \lfsr_c_0_a2_i_x2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[14]\, B => \tx_crc_data[0]\, C
         => N_161_i, D => N_228, Y => N_202_i_i);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \lfsr_c_0_a2_0_x2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[12]\, B => \tx_crc_data[11]\, C
         => N_520, D => N_519, Y => N_201_i);
    
    \lfsr_c_0_a2_2_x2[4]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[11]\, B => \tx_crc_data[10]\, C
         => N_519, D => N_518, Y => N_195_i);
    
    \lfsr_c_0_a2_1_0_x2[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => N_522, B => \tx_crc_data[15]\, Y => N_161_i);
    
    \lfsr_q[8]\ : SLE
      port map(D => N_202_i_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => N_9_0_i_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_crc_data[8]\);
    
    \lfsr_q[13]\ : SLE
      port map(D => \tx_crc_data[5]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => N_9_0_i_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_crc_data[13]\);
    
    \lfsr_c_0_a2[0]\ : CFG3
      generic map(INIT => x"96")

      port map(A => N_516, B => \lfsr_c[1]\, C => 
        \tx_crc_data[8]\, Y => \lfsr_c[0]\);
    
    \lfsr_q[15]\ : SLE
      port map(D => \lfsr_c[15]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => N_9_0_i_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_crc_data[15]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity TX_Collision_Detector is

    port( p2s_data              : in    std_logic_vector(7 downto 0);
          RX_FIFO_DIN           : in    std_logic_vector(7 downto 0);
          RX_FIFO_DIN_pipe_0    : in    std_logic;
          byte_clk_en_d_0       : in    std_logic;
          rx_crc_HighByte_en    : in    std_logic;
          DRVR_EN_c             : in    std_logic;
          N_6_0                 : in    std_logic;
          tx_col_detect_en      : out   std_logic;
          N_366_i               : in    std_logic;
          BIT_CLK               : in    std_logic;
          CommsFPGA_CCC_0_GL0   : in    std_logic;
          N_106_mux_i_i         : in    std_logic;
          TX_collision_detect_i : out   std_logic;
          TX_collision_detect   : out   std_logic
        );

end TX_Collision_Detector;

architecture DEF_ARCH of TX_Collision_Detector is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal TX_collision_detect_net_1, \RX_FIFO_wr_en_d[3]_net_1\, 
        VCC_net_1, \RX_FIFO_wr_en_d[2]_net_1\, GND_net_1, 
        \RX_FIFO_wr_en_d[4]_net_1\, \RX_FIFO_wr_en_d[5]_net_1\, 
        \RX_FIFO_wr_en_d[6]_net_1\, \RX_FIFO_wr_en_d[7]_net_1\, 
        \TX_FIFO_DOUT_d2_sync2RX[0]_net_1\, 
        \TX_FIFO_DOUT_d2[0]_net_1\, 
        \TX_FIFO_DOUT_d2_sync2RX[1]_net_1\, 
        \TX_FIFO_DOUT_d2[1]_net_1\, 
        \TX_FIFO_DOUT_d2_sync2RX[2]_net_1\, 
        \TX_FIFO_DOUT_d2[2]_net_1\, 
        \TX_FIFO_DOUT_d2_sync2RX[3]_net_1\, 
        \TX_FIFO_DOUT_d2[3]_net_1\, 
        \TX_FIFO_DOUT_d2_sync2RX[4]_net_1\, 
        \TX_FIFO_DOUT_d2[4]_net_1\, 
        \TX_FIFO_DOUT_d2_sync2RX[5]_net_1\, 
        \TX_FIFO_DOUT_d2[5]_net_1\, 
        \TX_FIFO_DOUT_d2_sync2RX[6]_net_1\, 
        \TX_FIFO_DOUT_d2[6]_net_1\, 
        \TX_FIFO_DOUT_d2_sync2RX[7]_net_1\, 
        \TX_FIFO_DOUT_d2[7]_net_1\, \TX_FIFO_DOUT_d1[6]_net_1\, 
        \TX_FIFO_DOUT_d1[7]_net_1\, \RX_FIFO_wr_en_d[0]_net_1\, 
        \RX_FIFO_wr_en_d[1]_net_1\, \RX_FIFO_DIN_d1[0]_net_1\, 
        \RX_FIFO_DIN_d1[1]_net_1\, \RX_FIFO_DIN_d1[2]_net_1\, 
        \RX_FIFO_DIN_d1[3]_net_1\, \RX_FIFO_DIN_d1[4]_net_1\, 
        \RX_FIFO_DIN_d1[5]_net_1\, \RX_FIFO_DIN_d1[6]_net_1\, 
        \RX_FIFO_DIN_d1[7]_net_1\, \TX_FIFO_DOUT_d1[0]_net_1\, 
        \TX_FIFO_DOUT_d1[1]_net_1\, \TX_FIFO_DOUT_d1[2]_net_1\, 
        \TX_FIFO_DOUT_d1[3]_net_1\, \TX_FIFO_DOUT_d1[4]_net_1\, 
        \TX_FIFO_DOUT_d1[5]_net_1\, 
        \TX_FIFO_DOUT_d2_syncCompare[0]_net_1\, 
        \TX_FIFO_DOUT_d2_syncCompare[1]_net_1\, 
        \TX_FIFO_DOUT_d2_syncCompare[2]_net_1\, 
        \TX_FIFO_DOUT_d2_syncCompare[3]_net_1\, 
        \TX_FIFO_DOUT_d2_syncCompare[4]_net_1\, 
        \TX_FIFO_DOUT_d2_syncCompare[5]_net_1\, 
        \TX_FIFO_DOUT_d2_syncCompare[6]_net_1\, 
        \TX_FIFO_DOUT_d2_syncCompare[7]_net_1\, 
        tx_collision_detect2, \un1_RX_FIFO_wr_en_d\, 
        \tx_col_detect_en_0\, un1_RX_FIFO_DIN_d1_NE_3, 
        un1_RX_FIFO_DIN_d1_NE_2, un1_RX_FIFO_DIN_d1_NE_1, 
        un1_RX_FIFO_DIN_d1_NE_0 : std_logic;

begin 

    TX_collision_detect <= TX_collision_detect_net_1;

    \RX_FIFO_DIN_d1[4]\ : SLE
      port map(D => RX_FIFO_DIN(4), CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_366_i, ALn => N_106_mux_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RX_FIFO_DIN_d1[4]_net_1\);
    
    \TX_FIFO_DOUT_d1[7]\ : SLE
      port map(D => p2s_data(7), CLK => BIT_CLK, EN => 
        byte_clk_en_d_0, ALn => N_106_mux_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \TX_FIFO_DOUT_d1[7]_net_1\);
    
    \RX_FIFO_wr_en_d[4]\ : SLE
      port map(D => \RX_FIFO_wr_en_d[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_wr_en_d[4]_net_1\);
    
    \RX_FIFO_wr_en_d[1]\ : SLE
      port map(D => \RX_FIFO_wr_en_d[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_wr_en_d[1]_net_1\);
    
    \RX_FIFO_wr_en_d[6]\ : SLE
      port map(D => \RX_FIFO_wr_en_d[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_wr_en_d[6]_net_1\);
    
    \TX_FIFO_DOUT_d2_syncCompare[1]\ : SLE
      port map(D => \TX_FIFO_DOUT_d2_sync2RX[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \RX_FIFO_wr_en_d[5]_net_1\, 
        ALn => N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_DOUT_d2_syncCompare[1]_net_1\);
    
    \TX_FIFO_DOUT_d2[2]\ : SLE
      port map(D => \TX_FIFO_DOUT_d1[2]_net_1\, CLK => BIT_CLK, 
        EN => byte_clk_en_d_0, ALn => N_106_mux_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \TX_FIFO_DOUT_d2[2]_net_1\);
    
    \TX_FIFO_DOUT_d1[2]\ : SLE
      port map(D => p2s_data(2), CLK => BIT_CLK, EN => 
        byte_clk_en_d_0, ALn => N_106_mux_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \TX_FIFO_DOUT_d1[2]_net_1\);
    
    \RX_FIFO_wr_en_d[2]\ : SLE
      port map(D => \RX_FIFO_wr_en_d[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_wr_en_d[2]_net_1\);
    
    \RX_FIFO_wr_en_d[5]\ : SLE
      port map(D => \RX_FIFO_wr_en_d[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_wr_en_d[5]_net_1\);
    
    \COLLISION_DETECT_PROC.un1_RX_FIFO_DIN_d1_NE_2\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => \TX_FIFO_DOUT_d2_syncCompare[5]_net_1\, B => 
        \TX_FIFO_DOUT_d2_syncCompare[4]_net_1\, C => 
        \RX_FIFO_DIN_d1[5]_net_1\, D => \RX_FIFO_DIN_d1[4]_net_1\, 
        Y => un1_RX_FIFO_DIN_d1_NE_2);
    
    \TX_FIFO_DOUT_d2_sync2RX[7]\ : SLE
      port map(D => \TX_FIFO_DOUT_d2[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_DOUT_d2_sync2RX[7]_net_1\);
    
    \RX_FIFO_DIN_d1[7]\ : SLE
      port map(D => RX_FIFO_DIN(7), CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_366_i, ALn => N_106_mux_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RX_FIFO_DIN_d1[7]_net_1\);
    
    \COLLISION_DETECT_PROC.un1_RX_FIFO_DIN_d1_NE\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => un1_RX_FIFO_DIN_d1_NE_3, B => 
        un1_RX_FIFO_DIN_d1_NE_2, C => un1_RX_FIFO_DIN_d1_NE_1, D
         => un1_RX_FIFO_DIN_d1_NE_0, Y => tx_collision_detect2);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \tx_col_detect_en\ : SLE
      port map(D => \tx_col_detect_en_0\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => tx_col_detect_en);
    
    TX_collision_detect_RNIAGUA : CFG1
      generic map(INIT => "01")

      port map(A => TX_collision_detect_net_1, Y => 
        TX_collision_detect_i);
    
    \TX_FIFO_DOUT_d1[5]\ : SLE
      port map(D => p2s_data(5), CLK => BIT_CLK, EN => 
        byte_clk_en_d_0, ALn => N_106_mux_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \TX_FIFO_DOUT_d1[5]_net_1\);
    
    \RX_FIFO_DIN_d1[1]\ : SLE
      port map(D => RX_FIFO_DIN(1), CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_366_i, ALn => N_106_mux_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RX_FIFO_DIN_d1[1]_net_1\);
    
    un1_RX_FIFO_wr_en_d : CFG3
      generic map(INIT => x"10")

      port map(A => rx_crc_HighByte_en, B => RX_FIFO_DIN_pipe_0, 
        C => \RX_FIFO_wr_en_d[7]_net_1\, Y => 
        \un1_RX_FIFO_wr_en_d\);
    
    \TX_FIFO_DOUT_d1[1]\ : SLE
      port map(D => p2s_data(1), CLK => BIT_CLK, EN => 
        byte_clk_en_d_0, ALn => N_106_mux_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \TX_FIFO_DOUT_d1[1]_net_1\);
    
    \RX_FIFO_DIN_d1[2]\ : SLE
      port map(D => RX_FIFO_DIN(2), CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_366_i, ALn => N_106_mux_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RX_FIFO_DIN_d1[2]_net_1\);
    
    \COLLISION_DETECT_PROC.un1_RX_FIFO_DIN_d1_NE_3\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => \TX_FIFO_DOUT_d2_syncCompare[7]_net_1\, B => 
        \TX_FIFO_DOUT_d2_syncCompare[6]_net_1\, C => 
        \RX_FIFO_DIN_d1[7]_net_1\, D => \RX_FIFO_DIN_d1[6]_net_1\, 
        Y => un1_RX_FIFO_DIN_d1_NE_3);
    
    \TX_FIFO_DOUT_d2_syncCompare[5]\ : SLE
      port map(D => \TX_FIFO_DOUT_d2_sync2RX[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \RX_FIFO_wr_en_d[5]_net_1\, 
        ALn => N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_DOUT_d2_syncCompare[5]_net_1\);
    
    \TX_FIFO_DOUT_d2_sync2RX[4]\ : SLE
      port map(D => \TX_FIFO_DOUT_d2[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_DOUT_d2_sync2RX[4]_net_1\);
    
    \TX_FIFO_DOUT_d2[0]\ : SLE
      port map(D => \TX_FIFO_DOUT_d1[0]_net_1\, CLK => BIT_CLK, 
        EN => byte_clk_en_d_0, ALn => N_106_mux_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \TX_FIFO_DOUT_d2[0]_net_1\);
    
    \TX_FIFO_DOUT_d2_syncCompare[7]\ : SLE
      port map(D => \TX_FIFO_DOUT_d2_sync2RX[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \RX_FIFO_wr_en_d[5]_net_1\, 
        ALn => N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_DOUT_d2_syncCompare[7]_net_1\);
    
    \TX_FIFO_DOUT_d2_sync2RX[1]\ : SLE
      port map(D => \TX_FIFO_DOUT_d2[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_DOUT_d2_sync2RX[1]_net_1\);
    
    \TX_FIFO_DOUT_d2[7]\ : SLE
      port map(D => \TX_FIFO_DOUT_d1[7]_net_1\, CLK => BIT_CLK, 
        EN => byte_clk_en_d_0, ALn => N_106_mux_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \TX_FIFO_DOUT_d2[7]_net_1\);
    
    tx_col_detect_en_0 : CFG2
      generic map(INIT => x"4")

      port map(A => N_6_0, B => DRVR_EN_c, Y => 
        \tx_col_detect_en_0\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \TX_FIFO_DOUT_d2_sync2RX[5]\ : SLE
      port map(D => \TX_FIFO_DOUT_d2[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_DOUT_d2_sync2RX[5]_net_1\);
    
    \TX_FIFO_DOUT_d2_syncCompare[4]\ : SLE
      port map(D => \TX_FIFO_DOUT_d2_sync2RX[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \RX_FIFO_wr_en_d[5]_net_1\, 
        ALn => N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_DOUT_d2_syncCompare[4]_net_1\);
    
    \TX_FIFO_DOUT_d2_syncCompare[0]\ : SLE
      port map(D => \TX_FIFO_DOUT_d2_sync2RX[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \RX_FIFO_wr_en_d[5]_net_1\, 
        ALn => N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_DOUT_d2_syncCompare[0]_net_1\);
    
    \RX_FIFO_wr_en_d[3]\ : SLE
      port map(D => \RX_FIFO_wr_en_d[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_wr_en_d[3]_net_1\);
    
    \TX_FIFO_DOUT_d2_syncCompare[2]\ : SLE
      port map(D => \TX_FIFO_DOUT_d2_sync2RX[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \RX_FIFO_wr_en_d[5]_net_1\, 
        ALn => N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_DOUT_d2_syncCompare[2]_net_1\);
    
    \RX_FIFO_DIN_d1[3]\ : SLE
      port map(D => RX_FIFO_DIN(3), CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_366_i, ALn => N_106_mux_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RX_FIFO_DIN_d1[3]_net_1\);
    
    \TX_FIFO_DOUT_d2[6]\ : SLE
      port map(D => \TX_FIFO_DOUT_d1[6]_net_1\, CLK => BIT_CLK, 
        EN => byte_clk_en_d_0, ALn => N_106_mux_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \TX_FIFO_DOUT_d2[6]_net_1\);
    
    \TX_FIFO_DOUT_d2_syncCompare[3]\ : SLE
      port map(D => \TX_FIFO_DOUT_d2_sync2RX[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \RX_FIFO_wr_en_d[5]_net_1\, 
        ALn => N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_DOUT_d2_syncCompare[3]_net_1\);
    
    \TX_FIFO_DOUT_d2[3]\ : SLE
      port map(D => \TX_FIFO_DOUT_d1[3]_net_1\, CLK => BIT_CLK, 
        EN => byte_clk_en_d_0, ALn => N_106_mux_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \TX_FIFO_DOUT_d2[3]_net_1\);
    
    \TX_FIFO_DOUT_d1[6]\ : SLE
      port map(D => p2s_data(6), CLK => BIT_CLK, EN => 
        byte_clk_en_d_0, ALn => N_106_mux_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \TX_FIFO_DOUT_d1[6]_net_1\);
    
    \RX_FIFO_wr_en_d[7]\ : SLE
      port map(D => \RX_FIFO_wr_en_d[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_wr_en_d[7]_net_1\);
    
    \RX_FIFO_DIN_d1[5]\ : SLE
      port map(D => RX_FIFO_DIN(5), CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_366_i, ALn => N_106_mux_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RX_FIFO_DIN_d1[5]_net_1\);
    
    \TX_collision_detect\ : SLE
      port map(D => tx_collision_detect2, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \un1_RX_FIFO_wr_en_d\, ALn => 
        N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        TX_collision_detect_net_1);
    
    \TX_FIFO_DOUT_d2[5]\ : SLE
      port map(D => \TX_FIFO_DOUT_d1[5]_net_1\, CLK => BIT_CLK, 
        EN => byte_clk_en_d_0, ALn => N_106_mux_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \TX_FIFO_DOUT_d2[5]_net_1\);
    
    \TX_FIFO_DOUT_d2[4]\ : SLE
      port map(D => \TX_FIFO_DOUT_d1[4]_net_1\, CLK => BIT_CLK, 
        EN => byte_clk_en_d_0, ALn => N_106_mux_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \TX_FIFO_DOUT_d2[4]_net_1\);
    
    \RX_FIFO_DIN_d1[6]\ : SLE
      port map(D => RX_FIFO_DIN(6), CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_366_i, ALn => N_106_mux_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RX_FIFO_DIN_d1[6]_net_1\);
    
    \TX_FIFO_DOUT_d2_sync2RX[2]\ : SLE
      port map(D => \TX_FIFO_DOUT_d2[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_DOUT_d2_sync2RX[2]_net_1\);
    
    \RX_FIFO_DIN_d1[0]\ : SLE
      port map(D => RX_FIFO_DIN(0), CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_366_i, ALn => N_106_mux_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RX_FIFO_DIN_d1[0]_net_1\);
    
    \COLLISION_DETECT_PROC.un1_RX_FIFO_DIN_d1_NE_0\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => \TX_FIFO_DOUT_d2_syncCompare[1]_net_1\, B => 
        \TX_FIFO_DOUT_d2_syncCompare[0]_net_1\, C => 
        \RX_FIFO_DIN_d1[1]_net_1\, D => \RX_FIFO_DIN_d1[0]_net_1\, 
        Y => un1_RX_FIFO_DIN_d1_NE_0);
    
    \TX_FIFO_DOUT_d2_sync2RX[3]\ : SLE
      port map(D => \TX_FIFO_DOUT_d2[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_DOUT_d2_sync2RX[3]_net_1\);
    
    \TX_FIFO_DOUT_d2_sync2RX[0]\ : SLE
      port map(D => \TX_FIFO_DOUT_d2[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_DOUT_d2_sync2RX[0]_net_1\);
    
    \COLLISION_DETECT_PROC.un1_RX_FIFO_DIN_d1_NE_1\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => \TX_FIFO_DOUT_d2_syncCompare[3]_net_1\, B => 
        \TX_FIFO_DOUT_d2_syncCompare[2]_net_1\, C => 
        \RX_FIFO_DIN_d1[3]_net_1\, D => \RX_FIFO_DIN_d1[2]_net_1\, 
        Y => un1_RX_FIFO_DIN_d1_NE_1);
    
    \TX_FIFO_DOUT_d1[3]\ : SLE
      port map(D => p2s_data(3), CLK => BIT_CLK, EN => 
        byte_clk_en_d_0, ALn => N_106_mux_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \TX_FIFO_DOUT_d1[3]_net_1\);
    
    \TX_FIFO_DOUT_d2[1]\ : SLE
      port map(D => \TX_FIFO_DOUT_d1[1]_net_1\, CLK => BIT_CLK, 
        EN => byte_clk_en_d_0, ALn => N_106_mux_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \TX_FIFO_DOUT_d2[1]_net_1\);
    
    \TX_FIFO_DOUT_d2_syncCompare[6]\ : SLE
      port map(D => \TX_FIFO_DOUT_d2_sync2RX[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \RX_FIFO_wr_en_d[5]_net_1\, 
        ALn => N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_DOUT_d2_syncCompare[6]_net_1\);
    
    \TX_FIFO_DOUT_d2_sync2RX[6]\ : SLE
      port map(D => \TX_FIFO_DOUT_d2[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        N_106_mux_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_DOUT_d2_sync2RX[6]_net_1\);
    
    \RX_FIFO_wr_en_d[0]\ : SLE
      port map(D => N_366_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => N_106_mux_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_wr_en_d[0]_net_1\);
    
    \TX_FIFO_DOUT_d1[4]\ : SLE
      port map(D => p2s_data(4), CLK => BIT_CLK, EN => 
        byte_clk_en_d_0, ALn => N_106_mux_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \TX_FIFO_DOUT_d1[4]_net_1\);
    
    \TX_FIFO_DOUT_d1[0]\ : SLE
      port map(D => p2s_data(0), CLK => BIT_CLK, EN => 
        byte_clk_en_d_0, ALn => N_106_mux_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \TX_FIFO_DOUT_d1[0]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity IdleLineDetectorZ0 is

    port( manches_in_dly      : in    std_logic_vector(1 downto 0);
          N_268_i             : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          N_480_i             : in    std_logic;
          tx_idle_line        : out   std_logic
        );

end IdleLineDetectorZ0;

architecture DEF_ARCH of IdleLineDetectorZ0 is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, N_339_i, GND_net_1, 
        \idle_line_cntr[0]_net_1\, \idle_line_cntr_s[0]\, 
        \idle_line_cntr[1]_net_1\, \idle_line_cntr_s[1]\, 
        \idle_line_cntr[2]_net_1\, \idle_line_cntr_s[2]\, 
        \idle_line_cntr[3]_net_1\, \idle_line_cntr_s[3]\, 
        \idle_line_cntr[4]_net_1\, \idle_line_cntr_s[4]\, 
        \idle_line_cntr[5]_net_1\, \idle_line_cntr_s[5]\, 
        \idle_line_cntr[6]_net_1\, \idle_line_cntr_s[6]_net_1\, 
        idle_line_cntr_cry_cy, \idle_line_cntr_cry_cy_Y[0]\, 
        un12_manches_in_dly, \N_268_i\, 
        \idle_line_cntr_cry[0]_net_1\, 
        \idle_line_cntr_cry[1]_net_1\, 
        \idle_line_cntr_cry[2]_net_1\, 
        \idle_line_cntr_cry[3]_net_1\, 
        \idle_line_cntr_cry[4]_net_1\, 
        \idle_line_cntr_cry[5]_net_1\, un12_manches_in_dly_4
         : std_logic;

begin 

    N_268_i <= \N_268_i\;

    idle_line_cntr_0_sqmuxa_i_x2 : CFG2
      generic map(INIT => x"6")

      port map(A => manches_in_dly(1), B => manches_in_dly(0), Y
         => \N_268_i\);
    
    \idle_line_cntr_cry[2]\ : ARI1
      generic map(INIT => x"4AC00")

      port map(A => VCC_net_1, B => \idle_line_cntr[2]_net_1\, C
         => N_339_i, D => \idle_line_cntr_cry_cy_Y[0]\, FCI => 
        \idle_line_cntr_cry[1]_net_1\, S => \idle_line_cntr_s[2]\, 
        Y => OPEN, FCO => \idle_line_cntr_cry[2]_net_1\);
    
    \idle_line_cntr[0]\ : SLE
      port map(D => \idle_line_cntr_s[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[0]_net_1\);
    
    idle_line : SLE
      port map(D => N_339_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        tx_idle_line);
    
    \idle_line_cntr_cry[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \idle_line_cntr[4]_net_1\, C
         => \idle_line_cntr_cry_cy_Y[0]\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[3]_net_1\, S => \idle_line_cntr_s[4]\, 
        Y => OPEN, FCO => \idle_line_cntr_cry[4]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \idle_line_cntr_cry[0]\ : ARI1
      generic map(INIT => x"48D88")

      port map(A => un12_manches_in_dly, B => 
        \idle_line_cntr_cry_cy_Y[0]\, C => 
        \idle_line_cntr[0]_net_1\, D => \N_268_i\, FCI => 
        idle_line_cntr_cry_cy, S => \idle_line_cntr_s[0]\, Y => 
        OPEN, FCO => \idle_line_cntr_cry[0]_net_1\);
    
    \idle_line_cntr_cry[3]\ : ARI1
      generic map(INIT => x"4AC00")

      port map(A => VCC_net_1, B => \idle_line_cntr[3]_net_1\, C
         => N_339_i, D => \idle_line_cntr_cry_cy_Y[0]\, FCI => 
        \idle_line_cntr_cry[2]_net_1\, S => \idle_line_cntr_s[3]\, 
        Y => OPEN, FCO => \idle_line_cntr_cry[3]_net_1\);
    
    \IDLE_LINE_DETECT_PROC.un12_manches_in_dly_RNI59RM\ : CFG2
      generic map(INIT => x"2")

      port map(A => un12_manches_in_dly, B => \N_268_i\, Y => 
        N_339_i);
    
    \idle_line_cntr_cry_cy[0]\ : ARI1
      generic map(INIT => x"41100")

      port map(A => VCC_net_1, B => un12_manches_in_dly, C => 
        \N_268_i\, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => \idle_line_cntr_cry_cy_Y[0]\, FCO => 
        idle_line_cntr_cry_cy);
    
    \idle_line_cntr_cry[1]\ : ARI1
      generic map(INIT => x"4AC00")

      port map(A => VCC_net_1, B => \idle_line_cntr[1]_net_1\, C
         => N_339_i, D => \idle_line_cntr_cry_cy_Y[0]\, FCI => 
        \idle_line_cntr_cry[0]_net_1\, S => \idle_line_cntr_s[1]\, 
        Y => OPEN, FCO => \idle_line_cntr_cry[1]_net_1\);
    
    \idle_line_cntr[4]\ : SLE
      port map(D => \idle_line_cntr_s[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[4]_net_1\);
    
    \IDLE_LINE_DETECT_PROC.un12_manches_in_dly\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \idle_line_cntr[6]_net_1\, B => 
        \idle_line_cntr[4]_net_1\, C => \idle_line_cntr[0]_net_1\, 
        D => un12_manches_in_dly_4, Y => un12_manches_in_dly);
    
    \idle_line_cntr_s[6]\ : ARI1
      generic map(INIT => x"4AC00")

      port map(A => VCC_net_1, B => \idle_line_cntr[6]_net_1\, C
         => N_339_i, D => \idle_line_cntr_cry_cy_Y[0]\, FCI => 
        \idle_line_cntr_cry[5]_net_1\, S => 
        \idle_line_cntr_s[6]_net_1\, Y => OPEN, FCO => OPEN);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \idle_line_cntr[6]\ : SLE
      port map(D => \idle_line_cntr_s[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[6]_net_1\);
    
    \idle_line_cntr[5]\ : SLE
      port map(D => \idle_line_cntr_s[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[5]_net_1\);
    
    \idle_line_cntr[1]\ : SLE
      port map(D => \idle_line_cntr_s[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[1]_net_1\);
    
    \idle_line_cntr[3]\ : SLE
      port map(D => \idle_line_cntr_s[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[3]_net_1\);
    
    \IDLE_LINE_DETECT_PROC.un12_manches_in_dly_4\ : CFG4
      generic map(INIT => x"4000")

      port map(A => \idle_line_cntr[5]_net_1\, B => 
        \idle_line_cntr[3]_net_1\, C => \idle_line_cntr[2]_net_1\, 
        D => \idle_line_cntr[1]_net_1\, Y => 
        un12_manches_in_dly_4);
    
    \idle_line_cntr_cry[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \idle_line_cntr[5]_net_1\, C
         => \idle_line_cntr_cry_cy_Y[0]\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[4]_net_1\, S => \idle_line_cntr_s[5]\, 
        Y => OPEN, FCO => \idle_line_cntr_cry[5]_net_1\);
    
    \idle_line_cntr[2]\ : SLE
      port map(D => \idle_line_cntr_s[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[2]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity TX_SM is

    port( manches_in_dly      : in    std_logic_vector(1 downto 0);
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          N_268_i             : out   std_logic;
          N_519               : in    std_logic;
          N_520               : in    std_logic;
          N_521               : in    std_logic;
          N_228               : in    std_logic;
          N_522               : in    std_logic;
          N_516               : in    std_logic;
          N_517               : in    std_logic;
          N_518               : in    std_logic;
          TX_FIFO_rd_en       : out   std_logic;
          TX_FIFO_Empty       : in    std_logic;
          TX_DataEn           : out   std_logic;
          TX_PreAmble         : out   std_logic;
          TX_PostAmble        : out   std_logic;
          tx_crc_byte1_en     : out   std_logic;
          tx_crc_byte2_en     : out   std_logic;
          tx_packet_complt    : out   std_logic;
          iTX_FIFO_rd_en      : out   std_logic;
          start_tx_FIFO       : in    std_logic;
          DRVR_EN_c           : out   std_logic;
          tx_crc_gen          : out   std_logic;
          byte_clk_en         : in    std_logic;
          tx_preamble_pat_en  : out   std_logic;
          BIT_CLK             : in    std_logic;
          N_480_i             : in    std_logic
        );

end TX_SM;

architecture DEF_ARCH of TX_SM is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IdleLineDetectorZ0
    port( manches_in_dly      : in    std_logic_vector(1 downto 0) := (others => 'U');
          N_268_i             : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          N_480_i             : in    std_logic := 'U';
          tx_idle_line        : out   std_logic
        );
  end component;

    signal \TX_STATE[8]_net_1\, \TX_STATE_i_0[8]\, 
        \PreAmble_cntr[1]_net_1\, VCC_net_1, N_132_i, GND_net_1, 
        \PreAmble_cntr[2]_net_1\, N_131_i, 
        \PreAmble_cntr[3]_net_1\, N_130_i, 
        \tx_packet_length[0]_net_1\, N_18_i, 
        un1_byte_clk_en_inv_2_i, \tx_packet_length[1]_net_1\, 
        N_22_i, \tx_packet_length[2]_net_1\, N_25_i, 
        \tx_packet_length[3]_net_1\, N_27_i, 
        \tx_packet_length[4]_net_1\, N_29_i, 
        \tx_packet_length[5]_net_1\, N_31_i, 
        \tx_packet_length[6]_net_1\, N_455_i, 
        \tx_packet_length[7]_net_1\, N_456_i, 
        \tx_packet_length[8]_net_1\, N_457_i, 
        \tx_packet_length[9]_net_1\, N_46_i, 
        \tx_packet_length[10]_net_1\, N_49_i, 
        \PostAmble_cntr[0]_net_1\, \PostAmble_cntr_34\, 
        \PostAmble_cntr[1]_net_1\, \PostAmble_cntr_35\, 
        \PostAmble_cntr[2]_net_1\, \PostAmble_cntr_36\, 
        \PreAmble_cntr[0]_net_1\, N_133_i, TX_DataEn_1_m, 
        \tx_byte_cntr_cry_cy_Y[0]\, \tx_idle_line_s\, 
        tx_idle_line, \start_tx_FIFO_s\, \TX_STATE[1]_net_1\, 
        \TX_STATE_62\, \TX_STATE[2]_net_1\, \TX_STATE_61\, 
        \TX_STATE[3]_net_1\, \TX_STATE_60\, \TX_STATE[4]_net_1\, 
        \TX_STATE_59\, \TX_STATE[5]_net_1\, \TX_STATE_58\, 
        \TX_STATE[6]_net_1\, \TX_STATE_57\, \TX_STATE[7]_net_1\, 
        \TX_STATE_56\, \TX_STATE_55\, iTX_FIFO_rd_en_net_1, 
        iTX_FIFO_rd_en_5, \TX_STATE[0]_net_1\, TX_DataEn_7, 
        \TX_STATE_63\, \tx_byte_cntr[0]_net_1\, 
        \tx_byte_cntr_s[0]\, \tx_byte_cntr[1]_net_1\, 
        \tx_byte_cntr_s[1]\, \tx_byte_cntr[2]_net_1\, 
        \tx_byte_cntr_s[2]\, \tx_byte_cntr[3]_net_1\, 
        \tx_byte_cntr_s[3]\, \tx_byte_cntr[4]_net_1\, 
        \tx_byte_cntr_s[4]\, \tx_byte_cntr[5]_net_1\, 
        \tx_byte_cntr_s[5]\, \tx_byte_cntr[6]_net_1\, 
        \tx_byte_cntr_s[6]\, \tx_byte_cntr[7]_net_1\, 
        \tx_byte_cntr_s[7]\, \tx_byte_cntr[8]_net_1\, 
        \tx_byte_cntr_s[8]\, \tx_byte_cntr[9]_net_1\, 
        \tx_byte_cntr_s[9]\, \tx_byte_cntr[10]_net_1\, 
        \tx_byte_cntr_s[10]\, \tx_byte_cntr[11]_net_1\, 
        \tx_byte_cntr_s[11]_net_1\, \txen_early_cntr[0]_net_1\, 
        \txen_early_cntr_s[0]\, \txen_early_cntr[1]_net_1\, 
        \txen_early_cntr_s[1]\, \txen_early_cntr[2]_net_1\, 
        \txen_early_cntr_s[2]\, \txen_early_cntr[3]_net_1\, 
        \txen_early_cntr_s[3]\, \txen_early_cntr[4]_net_1\, 
        \txen_early_cntr_s[4]\, \txen_early_cntr[5]_net_1\, 
        \txen_early_cntr_s[5]\, \txen_early_cntr[6]_net_1\, 
        \txen_early_cntr_s[6]\, \txen_early_cntr[7]_net_1\, 
        \txen_early_cntr_s[7]\, \txen_early_cntr[8]_net_1\, 
        \txen_early_cntr_s[8]\, \txen_early_cntr[9]_net_1\, 
        \txen_early_cntr_s[9]\, \txen_early_cntr[10]_net_1\, 
        \txen_early_cntr_s[10]\, \txen_early_cntr[11]_net_1\, 
        \txen_early_cntr_s[11]\, tx_byte_cntr_cry_cy, 
        \tx_byte_cntr_cry[0]_net_1\, \tx_byte_cntr_cry[1]_net_1\, 
        \tx_byte_cntr_cry[2]_net_1\, \tx_byte_cntr_cry[3]_net_1\, 
        \tx_byte_cntr_cry[4]_net_1\, \tx_byte_cntr_cry[5]_net_1\, 
        \tx_byte_cntr_cry[6]_net_1\, \tx_byte_cntr_cry[7]_net_1\, 
        \tx_byte_cntr_cry[8]_net_1\, \tx_byte_cntr_cry[9]_net_1\, 
        \tx_byte_cntr_cry[10]_net_1\, txen_early_cntr_cry_cy, 
        \TX_STATE_RNIAIGV2_Y[7]\, m15_e_6, m15_e_7, m15_e_8, 
        \txen_early_cntr_cry[0]\, \txen_early_cntr_cry[1]\, 
        \txen_early_cntr_cry[2]\, \txen_early_cntr_cry[3]\, 
        \txen_early_cntr_cry[4]\, \txen_early_cntr_cry[5]\, 
        \txen_early_cntr_cry[6]\, \txen_early_cntr_cry[7]\, 
        \txen_early_cntr_cry[8]\, \txen_early_cntr_cry[9]\, 
        \txen_early_cntr_cry[10]\, un26_tx_byte_cntr_a_4_cry_0, 
        un26_tx_byte_cntr_a_4_cry_1, \un26_tx_byte_cntr_a_4[2]\, 
        un26_tx_byte_cntr_a_4_cry_2, \un26_tx_byte_cntr_a_4[3]\, 
        un26_tx_byte_cntr_a_4_cry_3, \un26_tx_byte_cntr_a_4[4]\, 
        un26_tx_byte_cntr_a_4_cry_4, \un26_tx_byte_cntr_a_4[5]\, 
        un26_tx_byte_cntr_a_4_cry_5, \un26_tx_byte_cntr_a_4[6]\, 
        un26_tx_byte_cntr_a_4_cry_6, \un26_tx_byte_cntr_a_4[7]\, 
        un26_tx_byte_cntr_a_4_cry_7, \un26_tx_byte_cntr_a_4[8]\, 
        un26_tx_byte_cntr_a_4_cry_8, \un26_tx_byte_cntr_a_4[9]\, 
        un26_tx_byte_cntr_a_4_cry_9, \un26_tx_byte_cntr_a_4[10]\, 
        \un26_tx_byte_cntr_1_data_tmp[0]\, 
        \un26_tx_byte_cntr_1_data_tmp[1]\, 
        \un26_tx_byte_cntr_1_data_tmp[2]\, 
        \un26_tx_byte_cntr_1_data_tmp[3]\, N_235, 
        iTX_FIFO_rd_en_5_iv_0, N_93_i, N_13_i, un26_tx_byte_cntr, 
        \TX_STATE_58_1\, \TX_STATE_60_1\, N_568, 
        un10_tx_byte_cntr_0_a2_6_1, N_240, N_247, 
        un9_start_tx_fifo_s, N_252, N_484, N_489, 
        TX_STATE_3_sqmuxa, \un1_byte_clk_en_inv_2_0_2\, N_551, 
        N_161_i, un10_tx_byte_cntr_0_a2_5, N_552, N_232, 
        un15_tx_byte_cntr, N_454_i, un10_tx_byte_cntr, N_468_i, 
        N_464, un10_tx_byte_cntr_0_a2_6, N_487, N_256
         : std_logic;

    for all : IdleLineDetectorZ0
	Use entity work.IdleLineDetectorZ0(DEF_ARCH);
begin 

    iTX_FIFO_rd_en <= iTX_FIFO_rd_en_net_1;

    \TX_SM.un10_tx_byte_cntr_0_a2_6\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \tx_byte_cntr[11]_net_1\, B => 
        \tx_byte_cntr[8]_net_1\, C => \tx_byte_cntr[3]_net_1\, D
         => un10_tx_byte_cntr_0_a2_6_1, Y => 
        un10_tx_byte_cntr_0_a2_6);
    
    \TX_SM.un26_tx_byte_cntr_a_4_cry_5_RNIC95G3\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \tx_byte_cntr[7]_net_1\, B => 
        \un26_tx_byte_cntr_a_4[6]\, C => 
        \un26_tx_byte_cntr_a_4[7]\, D => \tx_byte_cntr[6]_net_1\, 
        FCI => \un26_tx_byte_cntr_1_data_tmp[2]\, S => OPEN, Y
         => OPEN, FCO => \un26_tx_byte_cntr_1_data_tmp[3]\);
    
    \tx_packet_length_RNO[2]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un15_tx_byte_cntr, B => N_518, C => 
        \tx_packet_length[2]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => N_25_i);
    
    \txen_early_cntr_RNIJFKLC[2]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[2]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[1]\, S => \txen_early_cntr_s[2]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[2]\);
    
    \PreAmble_cntr_RNO[0]\ : CFG4
      generic map(INIT => x"90AA")

      port map(A => \PreAmble_cntr[0]_net_1\, B => TX_FIFO_Empty, 
        C => \TX_STATE[6]_net_1\, D => byte_clk_en, Y => N_133_i);
    
    \tx_byte_cntr[8]\ : SLE
      port map(D => \tx_byte_cntr_s[8]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[8]_net_1\);
    
    \tx_byte_cntr[2]\ : SLE
      port map(D => \tx_byte_cntr_s[2]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[2]_net_1\);
    
    \TX_STATE[7]\ : SLE
      port map(D => \TX_STATE_56\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[7]_net_1\);
    
    \TX_SM.un26_tx_byte_cntr_a_4_cry_9\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \tx_packet_length[10]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        un26_tx_byte_cntr_a_4_cry_8, S => 
        \un26_tx_byte_cntr_a_4[10]\, Y => OPEN, FCO => 
        un26_tx_byte_cntr_a_4_cry_9);
    
    PostAmble_cntr_34 : CFG4
      generic map(INIT => x"04AA")

      port map(A => \PostAmble_cntr[0]_net_1\, B => 
        \TX_STATE[1]_net_1\, C => N_240, D => byte_clk_en, Y => 
        \PostAmble_cntr_34\);
    
    \TX_SM.PostAmble_cntr_9_i_o2[2]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \PostAmble_cntr[1]_net_1\, B => 
        \PostAmble_cntr[0]_net_1\, Y => N_489);
    
    \tx_byte_cntr_cry[7]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[7]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[6]_net_1\, S => \tx_byte_cntr_s[7]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[7]_net_1\);
    
    \TX_SM.un26_tx_byte_cntr_a_4_cry_0\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \tx_packet_length[1]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => GND_net_1, S => 
        OPEN, Y => OPEN, FCO => un26_tx_byte_cntr_a_4_cry_0);
    
    \PreAmble_cntr_RNO[2]\ : CFG4
      generic map(INIT => x"00A4")

      port map(A => \PreAmble_cntr[2]_net_1\, B => 
        \PreAmble_cntr[3]_net_1\, C => N_487, D => N_247, Y => 
        N_131_i);
    
    start_tx_FIFO_s : SLE
      port map(D => start_tx_FIFO, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \start_tx_FIFO_s\);
    
    \tx_packet_length[4]\ : SLE
      port map(D => N_29_i, CLK => BIT_CLK, EN => 
        un1_byte_clk_en_inv_2_i, ALn => N_480_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_packet_length[4]_net_1\);
    
    \tx_byte_cntr[0]\ : SLE
      port map(D => \tx_byte_cntr_s[0]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[0]_net_1\);
    
    \tx_packet_length[1]\ : SLE
      port map(D => N_22_i, CLK => BIT_CLK, EN => 
        un1_byte_clk_en_inv_2_i, ALn => N_480_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_packet_length[1]_net_1\);
    
    \TX_SM.un15_tx_byte_cntr_0_a5\ : CFG3
      generic map(INIT => x"80")

      port map(A => un10_tx_byte_cntr_0_a2_6, B => N_552, C => 
        un10_tx_byte_cntr_0_a2_5, Y => un15_tx_byte_cntr);
    
    \TX_SM.iTX_FIFO_rd_en_5_iv_1_0_0_a5\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_235, B => \TX_STATE[6]_net_1\, Y => 
        TX_DataEn_1_m);
    
    \txen_early_cntr_RNI5MOBM[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[5]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[4]\, S => \txen_early_cntr_s[5]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[5]\);
    
    un1_TX_STATE_7_i_a2_0_a5 : CFG4
      generic map(INIT => x"0001")

      port map(A => \TX_STATE[2]_net_1\, B => \TX_STATE[5]_net_1\, 
        C => \TX_STATE[4]_net_1\, D => \TX_STATE[3]_net_1\, Y => 
        N_161_i);
    
    \tx_byte_cntr_cry[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[4]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[3]_net_1\, S => \tx_byte_cntr_s[4]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[4]_net_1\);
    
    \TX_SM.iTX_FIFO_rd_en_5_iv\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => N_468_i, B => iTX_FIFO_rd_en_5_iv_0, C => 
        TX_STATE_3_sqmuxa, D => N_454_i, Y => iTX_FIFO_rd_en_5);
    
    \tx_packet_length_RNO[6]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un15_tx_byte_cntr, B => N_228, C => 
        \tx_packet_length[6]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => N_455_i);
    
    \un1_PreAmble_cntr_1_i_0_o2[1]\ : CFG3
      generic map(INIT => x"DF")

      port map(A => \PreAmble_cntr[1]_net_1\, B => N_484, C => 
        byte_clk_en, Y => N_487);
    
    \tx_packet_length_RNO[3]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un15_tx_byte_cntr, B => N_519, C => 
        \tx_packet_length[3]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => N_27_i);
    
    \TX_STATE[2]\ : SLE
      port map(D => \TX_STATE_61\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[2]_net_1\);
    
    \TX_PreAmble\ : SLE
      port map(D => \TX_STATE[6]_net_1\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        TX_PreAmble);
    
    \tx_packet_length[9]\ : SLE
      port map(D => N_46_i, CLK => BIT_CLK, EN => 
        un1_byte_clk_en_inv_2_i, ALn => N_480_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_packet_length[9]_net_1\);
    
    \txen_early_cntr_RNIFF8E9[1]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[1]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[0]\, S => \txen_early_cntr_s[1]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[1]\);
    
    \TX_SM.un26_tx_byte_cntr_a_4_cry_9_RNIP84Q\ : CFG4
      generic map(INIT => x"4812")

      port map(A => \tx_byte_cntr[11]_net_1\, B => 
        \tx_byte_cntr[10]_net_1\, C => 
        un26_tx_byte_cntr_a_4_cry_9, D => 
        \un26_tx_byte_cntr_a_4[10]\, Y => N_93_i);
    
    \txen_early_cntr[5]\ : SLE
      port map(D => \txen_early_cntr_s[5]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[5]_net_1\);
    
    TX_Enable : SLE
      port map(D => \TX_STATE_i_0[8]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        DRVR_EN_c);
    
    \tx_byte_cntr[6]\ : SLE
      port map(D => \tx_byte_cntr_s[6]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \tx_crc_byte2_en\ : SLE
      port map(D => \TX_STATE[2]_net_1\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        tx_crc_byte2_en);
    
    \tx_packet_length_RNO[0]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un15_tx_byte_cntr, B => N_516, C => 
        \tx_packet_length[0]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => N_18_i);
    
    \tx_byte_cntr_cry[10]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[10]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[9]_net_1\, S => \tx_byte_cntr_s[10]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[10]_net_1\);
    
    \tx_packet_length[3]\ : SLE
      port map(D => N_27_i, CLK => BIT_CLK, EN => 
        un1_byte_clk_en_inv_2_i, ALn => N_480_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_packet_length[3]_net_1\);
    
    \PreAmble_cntr[1]\ : SLE
      port map(D => N_132_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => N_480_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[1]_net_1\);
    
    \TX_SM.un26_tx_byte_cntr_a_4_cry_7\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \tx_packet_length[8]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        un26_tx_byte_cntr_a_4_cry_6, S => 
        \un26_tx_byte_cntr_a_4[8]\, Y => OPEN, FCO => 
        un26_tx_byte_cntr_a_4_cry_7);
    
    \TX_SM.PostAmble_cntr_9_i[1]\ : CFG4
      generic map(INIT => x"BF5F")

      port map(A => \PostAmble_cntr[0]_net_1\, B => 
        \PostAmble_cntr[2]_net_1\, C => \TX_STATE[1]_net_1\, D
         => \PostAmble_cntr[1]_net_1\, Y => N_464);
    
    \tx_byte_cntr_s[11]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[11]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[10]_net_1\, S => 
        \tx_byte_cntr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \iTX_FIFO_rd_en\ : SLE
      port map(D => iTX_FIFO_rd_en_5, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        iTX_FIFO_rd_en_net_1);
    
    \txen_early_cntr[8]\ : SLE
      port map(D => \txen_early_cntr_s[8]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[8]_net_1\);
    
    \tx_packet_length_RNO[1]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un15_tx_byte_cntr, B => N_517, C => 
        \tx_packet_length[1]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => N_22_i);
    
    \tx_byte_cntr[5]\ : SLE
      port map(D => \tx_byte_cntr_s[5]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[5]_net_1\);
    
    \TX_STATE[0]\ : SLE
      port map(D => \TX_STATE_63\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[0]_net_1\);
    
    \TX_SM.TX_DataEn_7_iv\ : CFG2
      generic map(INIT => x"B")

      port map(A => TX_DataEn_1_m, B => N_161_i, Y => TX_DataEn_7);
    
    \TX_STATE_ns_8_0_.m53_i_0_a2\ : CFG4
      generic map(INIT => x"E000")

      port map(A => N_551, B => N_552, C => 
        un10_tx_byte_cntr_0_a2_5, D => un10_tx_byte_cntr_0_a2_6, 
        Y => N_568);
    
    \tx_byte_cntr_cry[2]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[2]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[1]_net_1\, S => \tx_byte_cntr_s[2]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[2]_net_1\);
    
    \PreAmble_cntr[3]\ : SLE
      port map(D => N_130_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => N_480_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[3]_net_1\);
    
    \tx_packet_length[10]\ : SLE
      port map(D => N_49_i, CLK => BIT_CLK, EN => 
        un1_byte_clk_en_inv_2_i, ALn => N_480_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_packet_length[10]_net_1\);
    
    \txen_early_cntr_RNIUP0C61[10]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[10]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[9]\, S => \txen_early_cntr_s[10]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[10]\);
    
    \TX_SM.un26_tx_byte_cntr_a_4_cry_1_RNISDQP1\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \tx_byte_cntr[3]_net_1\, B => 
        \un26_tx_byte_cntr_a_4[2]\, C => 
        \un26_tx_byte_cntr_a_4[3]\, D => \tx_byte_cntr[2]_net_1\, 
        FCI => \un26_tx_byte_cntr_1_data_tmp[0]\, S => OPEN, Y
         => OPEN, FCO => \un26_tx_byte_cntr_1_data_tmp[1]\);
    
    \tx_byte_cntr[11]\ : SLE
      port map(D => \tx_byte_cntr_s[11]_net_1\, CLK => BIT_CLK, 
        EN => byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[11]_net_1\);
    
    \tx_byte_cntr_cry_cy[0]\ : ARI1
      generic map(INIT => x"4EE00")

      port map(A => VCC_net_1, B => \TX_STATE[4]_net_1\, C => 
        \TX_STATE[5]_net_1\, D => GND_net_1, FCI => VCC_net_1, S
         => OPEN, Y => \tx_byte_cntr_cry_cy_Y[0]\, FCO => 
        tx_byte_cntr_cry_cy);
    
    \tx_packet_length[5]\ : SLE
      port map(D => N_31_i, CLK => BIT_CLK, EN => 
        un1_byte_clk_en_inv_2_i, ALn => N_480_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_packet_length[5]_net_1\);
    
    \txen_early_cntr_RNIOG0TF[3]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[3]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[2]\, S => \txen_early_cntr_s[3]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[3]\);
    
    TX_STATE_58 : CFG4
      generic map(INIT => x"4CEE")

      port map(A => byte_clk_en, B => \TX_STATE[5]_net_1\, C => 
        un26_tx_byte_cntr, D => \TX_STATE_58_1\, Y => 
        \TX_STATE_58\);
    
    TX_STATE_58_1 : CFG3
      generic map(INIT => x"15")

      port map(A => \TX_STATE[4]_net_1\, B => \TX_STATE[5]_net_1\, 
        C => N_568, Y => \TX_STATE_58_1\);
    
    \txen_early_cntr[9]\ : SLE
      port map(D => \txen_early_cntr_s[9]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[9]_net_1\);
    
    \TX_STATE_RNIAIGV2[7]\ : ARI1
      generic map(INIT => x"42AAA")

      port map(A => m15_e_8, B => \TX_STATE[7]_net_1\, C => 
        m15_e_6, D => m15_e_7, FCI => VCC_net_1, S => OPEN, Y => 
        \TX_STATE_RNIAIGV2_Y[7]\, FCO => txen_early_cntr_cry_cy);
    
    TX_STATE_60_1 : CFG2
      generic map(INIT => x"4")

      port map(A => N_568, B => \TX_STATE[5]_net_1\, Y => 
        \TX_STATE_60_1\);
    
    \PreAmble_cntr_RNO[3]\ : CFG4
      generic map(INIT => x"00C6")

      port map(A => \PreAmble_cntr[2]_net_1\, B => 
        \PreAmble_cntr[3]_net_1\, C => N_487, D => N_247, Y => 
        N_130_i);
    
    \TX_STATE_ns_8_0_.m59_i_o2\ : CFG3
      generic map(INIT => x"FD")

      port map(A => \PostAmble_cntr[1]_net_1\, B => 
        \PostAmble_cntr[2]_net_1\, C => \PostAmble_cntr[0]_net_1\, 
        Y => N_232);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \tx_byte_cntr[4]\ : SLE
      port map(D => \tx_byte_cntr_s[4]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[4]_net_1\);
    
    \TX_SM.iTX_FIFO_rd_en_5_iv_RNO\ : CFG2
      generic map(INIT => x"8")

      port map(A => un10_tx_byte_cntr, B => \TX_STATE[5]_net_1\, 
        Y => N_468_i);
    
    \txen_early_cntr[1]\ : SLE
      port map(D => \txen_early_cntr_s[1]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[1]_net_1\);
    
    \tx_byte_cntr_cry[0]\ : ARI1
      generic map(INIT => x"4A800")

      port map(A => VCC_net_1, B => \tx_byte_cntr[0]_net_1\, C
         => \TX_STATE[5]_net_1\, D => \TX_STATE[4]_net_1\, FCI
         => tx_byte_cntr_cry_cy, S => \tx_byte_cntr_s[0]\, Y => 
        OPEN, FCO => \tx_byte_cntr_cry[0]_net_1\);
    
    \TX_STATE_ns_8_0_.m15_e_6\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \txen_early_cntr[5]_net_1\, B => 
        \txen_early_cntr[4]_net_1\, C => 
        \txen_early_cntr[3]_net_1\, D => 
        \txen_early_cntr[2]_net_1\, Y => m15_e_6);
    
    \txen_early_cntr_RNIBD9931[9]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[9]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[8]\, S => \txen_early_cntr_s[9]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[9]\);
    
    \tx_packet_length[8]\ : SLE
      port map(D => N_457_i, CLK => BIT_CLK, EN => 
        un1_byte_clk_en_inv_2_i, ALn => N_480_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_packet_length[8]_net_1\);
    
    \tx_byte_cntr_cry[1]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[1]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[0]_net_1\, S => \tx_byte_cntr_s[1]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[1]_net_1\);
    
    \TX_SM.un26_tx_byte_cntr_a_4_cry_4\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \tx_packet_length[5]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        un26_tx_byte_cntr_a_4_cry_3, S => 
        \un26_tx_byte_cntr_a_4[5]\, Y => OPEN, FCO => 
        un26_tx_byte_cntr_a_4_cry_4);
    
    \TX_DataEn\ : SLE
      port map(D => TX_DataEn_7, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        TX_DataEn);
    
    \tx_byte_cntr[3]\ : SLE
      port map(D => \tx_byte_cntr_s[3]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[3]_net_1\);
    
    \tx_byte_cntr[7]\ : SLE
      port map(D => \tx_byte_cntr_s[7]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[7]_net_1\);
    
    \TX_SM.un10_tx_byte_cntr_0_a5\ : CFG3
      generic map(INIT => x"80")

      port map(A => un10_tx_byte_cntr_0_a2_6, B => N_551, C => 
        un10_tx_byte_cntr_0_a2_5, Y => un10_tx_byte_cntr);
    
    \TX_SM.un26_tx_byte_cntr_a_4_cry_7_RNI4K5R\ : CFG4
      generic map(INIT => x"8241")

      port map(A => \tx_byte_cntr[8]_net_1\, B => 
        \tx_byte_cntr[9]_net_1\, C => \un26_tx_byte_cntr_a_4[9]\, 
        D => \un26_tx_byte_cntr_a_4[8]\, Y => N_13_i);
    
    TX_STATE_61 : CFG3
      generic map(INIT => x"E2")

      port map(A => \TX_STATE[2]_net_1\, B => byte_clk_en, C => 
        \TX_STATE[3]_net_1\, Y => \TX_STATE_61\);
    
    \TX_STATE[8]\ : SLE
      port map(D => \TX_STATE_55\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[8]_net_1\);
    
    \txen_early_cntr_RNIDQ4JP[6]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[6]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[5]\, S => \txen_early_cntr_s[6]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[6]\);
    
    \txen_early_cntr_RNO[11]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[11]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[10]\, S => \txen_early_cntr_s[11]\, 
        Y => OPEN, FCO => OPEN);
    
    \txen_early_cntr_RNICGS66[0]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[0]_net_1\, D => GND_net_1, FCI => 
        txen_early_cntr_cry_cy, S => \txen_early_cntr_s[0]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[0]\);
    
    \tx_packet_complt\ : SLE
      port map(D => \TX_STATE[0]_net_1\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        tx_packet_complt);
    
    TX_STATE_55 : CFG4
      generic map(INIT => x"FC70")

      port map(A => un9_start_tx_fifo_s, B => byte_clk_en, C => 
        \TX_STATE[8]_net_1\, D => \TX_STATE[0]_net_1\, Y => 
        \TX_STATE_55\);
    
    \txen_early_cntr[0]\ : SLE
      port map(D => \txen_early_cntr_s[0]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[0]_net_1\);
    
    \TX_SM.un26_tx_byte_cntr_a_4_cry_6\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \tx_packet_length[7]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        un26_tx_byte_cntr_a_4_cry_5, S => 
        \un26_tx_byte_cntr_a_4[7]\, Y => OPEN, FCO => 
        un26_tx_byte_cntr_a_4_cry_6);
    
    PostAmble_cntr_35 : CFG3
      generic map(INIT => x"5C")

      port map(A => N_464, B => \PostAmble_cntr[1]_net_1\, C => 
        byte_clk_en, Y => \PostAmble_cntr_35\);
    
    \TX_STATE_ns_8_0_.m15_e_7\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \txen_early_cntr[11]_net_1\, B => 
        \txen_early_cntr[10]_net_1\, C => 
        \txen_early_cntr[1]_net_1\, D => 
        \txen_early_cntr[0]_net_1\, Y => m15_e_7);
    
    \PreAmble_cntr[2]\ : SLE
      port map(D => N_131_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => N_480_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[2]_net_1\);
    
    TX_STATE_62 : CFG4
      generic map(INIT => x"EACA")

      port map(A => \TX_STATE[1]_net_1\, B => \TX_STATE[2]_net_1\, 
        C => byte_clk_en, D => N_232, Y => \TX_STATE_62\);
    
    \TX_STATE_ns_8_0_.m16_i_0_a5_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => un9_start_tx_fifo_s, B => \TX_STATE[8]_net_1\, 
        Y => N_252);
    
    \TX_STATE_ns_8_0_.m51_i_0_a5_0\ : CFG2
      generic map(INIT => x"4")

      port map(A => un26_tx_byte_cntr, B => \TX_STATE[5]_net_1\, 
        Y => TX_STATE_3_sqmuxa);
    
    \un1_PreAmble_cntr_1_i_0_a5_0[1]\ : CFG2
      generic map(INIT => x"2")

      port map(A => byte_clk_en, B => \TX_STATE[6]_net_1\, Y => 
        N_247);
    
    \TX_SM.iTX_FIFO_rd_en_5_iv_0\ : CFG3
      generic map(INIT => x"DC")

      port map(A => N_235, B => \TX_STATE[4]_net_1\, C => 
        \TX_STATE[6]_net_1\, Y => iTX_FIFO_rd_en_5_iv_0);
    
    \tx_packet_length[6]\ : SLE
      port map(D => N_455_i, CLK => BIT_CLK, EN => 
        un1_byte_clk_en_inv_2_i, ALn => N_480_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_packet_length[6]_net_1\);
    
    \tx_byte_cntr[10]\ : SLE
      port map(D => \tx_byte_cntr_s[10]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[10]_net_1\);
    
    \TX_SM.un26_tx_byte_cntr_a_4_cry_3_RNIGPVK2\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \tx_byte_cntr[5]_net_1\, B => 
        \un26_tx_byte_cntr_a_4[4]\, C => 
        \un26_tx_byte_cntr_a_4[5]\, D => \tx_byte_cntr[4]_net_1\, 
        FCI => \un26_tx_byte_cntr_1_data_tmp[1]\, S => OPEN, Y
         => OPEN, FCO => \un26_tx_byte_cntr_1_data_tmp[2]\);
    
    PostAmble_cntr_36 : CFG4
      generic map(INIT => x"84AA")

      port map(A => \PostAmble_cntr[2]_net_1\, B => 
        \TX_STATE[1]_net_1\, C => N_489, D => byte_clk_en, Y => 
        \PostAmble_cntr_36\);
    
    un1_byte_clk_en_inv_2_0_2 : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \TX_STATE[2]_net_1\, B => byte_clk_en, C => 
        \TX_STATE[4]_net_1\, D => \TX_STATE[3]_net_1\, Y => 
        \un1_byte_clk_en_inv_2_0_2\);
    
    un1_byte_clk_en_inv_2_0_2_RNIJ5S61 : CFG4
      generic map(INIT => x"3331")

      port map(A => \TX_STATE[5]_net_1\, B => 
        \un1_byte_clk_en_inv_2_0_2\, C => un10_tx_byte_cntr, D
         => un15_tx_byte_cntr, Y => un1_byte_clk_en_inv_2_i);
    
    \TX_STATE_ns_8_0_.m15_e_8\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \txen_early_cntr[9]_net_1\, B => 
        \txen_early_cntr[8]_net_1\, C => 
        \txen_early_cntr[7]_net_1\, D => 
        \txen_early_cntr[6]_net_1\, Y => m15_e_8);
    
    \TX_SM.un26_tx_byte_cntr_a_4_cry_8\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \tx_packet_length[9]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        un26_tx_byte_cntr_a_4_cry_7, S => 
        \un26_tx_byte_cntr_a_4[9]\, Y => OPEN, FCO => 
        un26_tx_byte_cntr_a_4_cry_8);
    
    \TX_SM.un26_tx_byte_cntr_a_4_cry_1\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \tx_packet_length[2]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        un26_tx_byte_cntr_a_4_cry_0, S => 
        \un26_tx_byte_cntr_a_4[2]\, Y => OPEN, FCO => 
        un26_tx_byte_cntr_a_4_cry_1);
    
    TX_STATE_57 : CFG4
      generic map(INIT => x"EAF0")

      port map(A => N_256, B => N_235, C => \TX_STATE[6]_net_1\, 
        D => byte_clk_en, Y => \TX_STATE_57\);
    
    \txen_early_cntr[4]\ : SLE
      port map(D => \txen_early_cntr_s[4]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[4]_net_1\);
    
    \tx_crc_byte1_en\ : SLE
      port map(D => \TX_STATE[3]_net_1\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        tx_crc_byte1_en);
    
    \tx_byte_cntr_cry[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[5]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[4]_net_1\, S => \tx_byte_cntr_s[5]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[5]_net_1\);
    
    \PostAmble_cntr[2]\ : SLE
      port map(D => \PostAmble_cntr_36\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PostAmble_cntr[2]_net_1\);
    
    TX_STATE_56 : CFG4
      generic map(INIT => x"EEF0")

      port map(A => N_252, B => \TX_STATE_RNIAIGV2_Y[7]\, C => 
        \TX_STATE[7]_net_1\, D => byte_clk_en, Y => \TX_STATE_56\);
    
    \PostAmble_cntr[1]\ : SLE
      port map(D => \PostAmble_cntr_35\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PostAmble_cntr[1]_net_1\);
    
    \txen_early_cntr[2]\ : SLE
      port map(D => \txen_early_cntr_s[2]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[2]_net_1\);
    
    TX_STATE_60 : CFG4
      generic map(INIT => x"E444")

      port map(A => byte_clk_en, B => \TX_STATE[3]_net_1\, C => 
        un26_tx_byte_cntr, D => \TX_STATE_60_1\, Y => 
        \TX_STATE_60\);
    
    \TX_SM.un15_tx_byte_cntr_0_a5_0\ : CFG3
      generic map(INIT => x"02")

      port map(A => \tx_byte_cntr[2]_net_1\, B => 
        \tx_byte_cntr[1]_net_1\, C => \tx_byte_cntr[0]_net_1\, Y
         => N_552);
    
    \tx_packet_length[2]\ : SLE
      port map(D => N_25_i, CLK => BIT_CLK, EN => 
        un1_byte_clk_en_inv_2_i, ALn => N_480_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_packet_length[2]_net_1\);
    
    \txen_early_cntr_RNIUIC4J[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[4]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[3]\, S => \txen_early_cntr_s[4]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[4]\);
    
    \tx_byte_cntr_cry[6]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[6]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[5]_net_1\, S => \tx_byte_cntr_s[6]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[6]_net_1\);
    
    \un1_PreAmble_cntr_1_i_0_o2_0[0]\ : CFG2
      generic map(INIT => x"B")

      port map(A => TX_FIFO_Empty, B => \PreAmble_cntr[0]_net_1\, 
        Y => N_484);
    
    \txen_early_cntr[7]\ : SLE
      port map(D => \txen_early_cntr_s[7]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[7]_net_1\);
    
    \txen_early_cntr[3]\ : SLE
      port map(D => \txen_early_cntr_s[3]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[3]_net_1\);
    
    \tx_packet_length_RNO[8]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un15_tx_byte_cntr, B => N_516, C => 
        \tx_packet_length[8]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => N_457_i);
    
    \TX_SM.un26_tx_byte_cntr_a_4_cry_5_RNI96F55\ : CFG3
      generic map(INIT => x"20")

      port map(A => N_93_i, B => 
        \un26_tx_byte_cntr_1_data_tmp[3]\, C => N_13_i, Y => 
        un26_tx_byte_cntr);
    
    iTX_PostAmble : SLE
      port map(D => \TX_STATE[1]_net_1\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        TX_PostAmble);
    
    TX_STATE_63 : CFG4
      generic map(INIT => x"0CAA")

      port map(A => \TX_STATE[0]_net_1\, B => \TX_STATE[1]_net_1\, 
        C => N_232, D => byte_clk_en, Y => \TX_STATE_63\);
    
    \tx_packet_length_RNO[5]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un15_tx_byte_cntr, B => N_521, C => 
        \tx_packet_length[5]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => N_31_i);
    
    \tx_packet_length_RNO[7]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un15_tx_byte_cntr, B => N_522, C => 
        \tx_packet_length[7]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => N_456_i);
    
    \tx_packet_length_RNO[9]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un15_tx_byte_cntr, B => N_517, C => 
        \tx_packet_length[9]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => N_46_i);
    
    \tx_byte_cntr[1]\ : SLE
      port map(D => \tx_byte_cntr_s[1]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[1]_net_1\);
    
    \TX_SM.un10_tx_byte_cntr_0_a2_5\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \tx_byte_cntr[7]_net_1\, B => 
        \tx_byte_cntr[6]_net_1\, C => \tx_byte_cntr[5]_net_1\, D
         => \tx_byte_cntr[4]_net_1\, Y => 
        un10_tx_byte_cntr_0_a2_5);
    
    \txen_early_cntr_RNI06T101[8]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[8]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[7]\, S => \txen_early_cntr_s[8]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[8]\);
    
    \PreAmble_cntr[0]\ : SLE
      port map(D => N_133_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => N_480_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[0]_net_1\);
    
    \PostAmble_cntr[0]\ : SLE
      port map(D => \PostAmble_cntr_34\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PostAmble_cntr[0]_net_1\);
    
    \TX_SM.un26_tx_byte_cntr_a_4_cry_2\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \tx_packet_length[3]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        un26_tx_byte_cntr_a_4_cry_1, S => 
        \un26_tx_byte_cntr_a_4[3]\, Y => OPEN, FCO => 
        un26_tx_byte_cntr_a_4_cry_2);
    
    \tx_crc_gen\ : SLE
      port map(D => \tx_byte_cntr_cry_cy_Y[0]\, CLK => BIT_CLK, 
        EN => byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        tx_crc_gen);
    
    \TX_STATE_ns_8_0_.m53_i_0_a2_0\ : CFG3
      generic map(INIT => x"40")

      port map(A => \tx_byte_cntr[2]_net_1\, B => 
        \tx_byte_cntr[1]_net_1\, C => \tx_byte_cntr[0]_net_1\, Y
         => N_551);
    
    \TX_STATE[4]\ : SLE
      port map(D => \TX_STATE_59\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[4]_net_1\);
    
    \tx_packet_length[7]\ : SLE
      port map(D => N_456_i, CLK => BIT_CLK, EN => 
        un1_byte_clk_en_inv_2_i, ALn => N_480_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_packet_length[7]_net_1\);
    
    \TX_STATE[5]\ : SLE
      port map(D => \TX_STATE_58\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[5]_net_1\);
    
    \tx_packet_length_RNO[4]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => un15_tx_byte_cntr, B => N_520, C => 
        \tx_packet_length[4]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => N_29_i);
    
    \txen_early_cntr[10]\ : SLE
      port map(D => \txen_early_cntr_s[10]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[10]_net_1\);
    
    \TX_STATE[3]\ : SLE
      port map(D => \TX_STATE_60\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[3]_net_1\);
    
    \tx_packet_length_RNO[10]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => un15_tx_byte_cntr, B => N_518, C => 
        \tx_packet_length[10]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => N_49_i);
    
    \tx_byte_cntr_cry[9]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[9]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[8]_net_1\, S => \tx_byte_cntr_s[9]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[9]_net_1\);
    
    \PreAmble_cntr_RNO[1]\ : CFG4
      generic map(INIT => x"090C")

      port map(A => N_484, B => \PreAmble_cntr[1]_net_1\, C => 
        N_247, D => byte_clk_en, Y => N_132_i);
    
    \TX_SM.un26_tx_byte_cntr_a_4_cry_3\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \tx_packet_length[4]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        un26_tx_byte_cntr_a_4_cry_2, S => 
        \un26_tx_byte_cntr_a_4[4]\, Y => OPEN, FCO => 
        un26_tx_byte_cntr_a_4_cry_3);
    
    TX_Enable_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \TX_STATE[8]_net_1\, Y => \TX_STATE_i_0[8]\);
    
    \tx_packet_length_RNIG6LU[0]\ : ARI1
      generic map(INIT => x"62184")

      port map(A => \tx_packet_length[1]_net_1\, B => 
        \tx_byte_cntr[0]_net_1\, C => \tx_byte_cntr[1]_net_1\, D
         => \tx_packet_length[0]_net_1\, FCI => GND_net_1, S => 
        OPEN, Y => OPEN, FCO => \un26_tx_byte_cntr_1_data_tmp[0]\);
    
    TX_IDLE_LINE_DETECTOR : IdleLineDetectorZ0
      port map(manches_in_dly(1) => manches_in_dly(1), 
        manches_in_dly(0) => manches_in_dly(0), N_268_i => 
        N_268_i, CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        N_480_i => N_480_i, tx_idle_line => tx_idle_line);
    
    tx_idle_line_s : SLE
      port map(D => tx_idle_line, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_idle_line_s\);
    
    \TX_SM.PostAmble_cntr_9_i_a5[0]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \PostAmble_cntr[1]_net_1\, B => 
        \PostAmble_cntr[2]_net_1\, Y => N_240);
    
    \tx_packet_length[0]\ : SLE
      port map(D => N_18_i, CLK => BIT_CLK, EN => 
        un1_byte_clk_en_inv_2_i, ALn => N_480_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_packet_length[0]_net_1\);
    
    \TX_SM.un9_start_tx_fifo_s\ : CFG2
      generic map(INIT => x"8")

      port map(A => \start_tx_FIFO_s\, B => \tx_idle_line_s\, Y
         => un9_start_tx_fifo_s);
    
    \txen_early_cntr[6]\ : SLE
      port map(D => \txen_early_cntr_s[6]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[6]_net_1\);
    
    \TX_SM.un26_tx_byte_cntr_a_4_cry_5\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \tx_packet_length[6]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        un26_tx_byte_cntr_a_4_cry_4, S => 
        \un26_tx_byte_cntr_a_4[6]\, Y => OPEN, FCO => 
        un26_tx_byte_cntr_a_4_cry_5);
    
    \tx_byte_cntr[9]\ : SLE
      port map(D => \tx_byte_cntr_s[9]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[9]_net_1\);
    
    \tx_byte_cntr_cry[8]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[8]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[7]_net_1\, S => \tx_byte_cntr_s[8]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[8]_net_1\);
    
    \tx_byte_cntr_cry[3]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[3]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[2]_net_1\, S => \tx_byte_cntr_s[3]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[3]_net_1\);
    
    \TX_SM.un10_tx_byte_cntr_0_a2_6_1\ : CFG2
      generic map(INIT => x"1")

      port map(A => \tx_byte_cntr[9]_net_1\, B => 
        \tx_byte_cntr[10]_net_1\, Y => un10_tx_byte_cntr_0_a2_6_1);
    
    \txen_early_cntr_RNIMVGQS[7]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[7]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[6]\, S => \txen_early_cntr_s[7]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[7]\);
    
    \TX_STATE_ns_8_0_.m35_i_0_o2\ : CFG4
      generic map(INIT => x"FFFD")

      port map(A => \PreAmble_cntr[1]_net_1\, B => N_484, C => 
        \PreAmble_cntr[3]_net_1\, D => \PreAmble_cntr[2]_net_1\, 
        Y => N_235);
    
    \TX_STATE_ns_8_0_.m35_i_0_a5_0\ : CFG4
      generic map(INIT => x"8000")

      port map(A => m15_e_7, B => m15_e_6, C => 
        \TX_STATE[7]_net_1\, D => m15_e_8, Y => N_256);
    
    \TX_STATE[6]\ : SLE
      port map(D => \TX_STATE_57\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[6]_net_1\);
    
    \tx_preamble_pat_en\ : SLE
      port map(D => TX_DataEn_1_m, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        tx_preamble_pat_en);
    
    \TX_STATE[1]\ : SLE
      port map(D => \TX_STATE_62\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[1]_net_1\);
    
    TX_STATE_59 : CFG3
      generic map(INIT => x"D8")

      port map(A => byte_clk_en, B => TX_DataEn_1_m, C => 
        \TX_STATE[4]_net_1\, Y => \TX_STATE_59\);
    
    \TX_SM.iTX_FIFO_rd_en_5_iv_RNO_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => un15_tx_byte_cntr, B => \TX_STATE[5]_net_1\, 
        Y => N_454_i);
    
    \txen_early_cntr[11]\ : SLE
      port map(D => \txen_early_cntr_s[11]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => N_480_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[11]_net_1\);
    
    \TX_FIFO_rd_en\ : CFG2
      generic map(INIT => x"8")

      port map(A => byte_clk_en, B => iTX_FIFO_rd_en_net_1, Y => 
        TX_FIFO_rd_en);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity ManchesEncoder is

    port( manches_in_dly        : in    std_logic_vector(1 downto 0);
          RX_FIFO_DIN           : in    std_logic_vector(7 downto 0);
          RX_FIFO_DIN_pipe_0    : in    std_logic;
          p2s_data_0            : out   std_logic;
          N_9_0_i_i             : in    std_logic;
          start_tx_FIFO         : in    std_logic;
          iTX_FIFO_rd_en        : out   std_logic;
          tx_packet_complt      : out   std_logic;
          TX_PreAmble           : out   std_logic;
          TX_FIFO_Empty         : in    std_logic;
          TX_FIFO_rd_en         : out   std_logic;
          N_268_i               : out   std_logic;
          TX_collision_detect   : out   std_logic;
          TX_collision_detect_i : out   std_logic;
          N_106_mux_i_i         : in    std_logic;
          CommsFPGA_CCC_0_GL0   : in    std_logic;
          N_366_i               : in    std_logic;
          tx_col_detect_en      : out   std_logic;
          N_6_0                 : in    std_logic;
          DRVR_EN_c             : out   std_logic;
          rx_crc_HighByte_en    : in    std_logic;
          un19_tx_dataen        : out   std_logic;
          N_517                 : in    std_logic;
          N_522                 : in    std_logic;
          N_519                 : in    std_logic;
          N_518                 : in    std_logic;
          N_521                 : in    std_logic;
          N_520                 : in    std_logic;
          N_228                 : in    std_logic;
          N_516                 : in    std_logic;
          tx_preamble_pat_en    : out   std_logic;
          TX_PostAmble_d1       : out   std_logic;
          MANCHESTER_OUT_5      : in    std_logic;
          CommsFPGA_CCC_0_GL1   : in    std_logic;
          byte_clk_en           : in    std_logic;
          BIT_CLK               : in    std_logic;
          N_480_i               : in    std_logic;
          MANCH_OUT_P_c_i       : out   std_logic;
          MANCH_OUT_P_c         : out   std_logic
        );

end ManchesEncoder;

architecture DEF_ARCH of ManchesEncoder is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CRC16_Generator_0
    port( tx_crc_data : out   std_logic_vector(15 downto 0);
          N_518       : in    std_logic := 'U';
          N_519       : in    std_logic := 'U';
          N_228       : in    std_logic := 'U';
          N_520       : in    std_logic := 'U';
          N_521       : in    std_logic := 'U';
          N_516       : in    std_logic := 'U';
          N_517       : in    std_logic := 'U';
          N_522       : in    std_logic := 'U';
          tx_crc_gen  : in    std_logic := 'U';
          byte_clk_en : in    std_logic := 'U';
          BIT_CLK     : in    std_logic := 'U';
          N_9_0_i_i   : in    std_logic := 'U'
        );
  end component;

  component TX_Collision_Detector
    port( p2s_data              : in    std_logic_vector(7 downto 0) := (others => 'U');
          RX_FIFO_DIN           : in    std_logic_vector(7 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe_0    : in    std_logic := 'U';
          byte_clk_en_d_0       : in    std_logic := 'U';
          rx_crc_HighByte_en    : in    std_logic := 'U';
          DRVR_EN_c             : in    std_logic := 'U';
          N_6_0                 : in    std_logic := 'U';
          tx_col_detect_en      : out   std_logic;
          N_366_i               : in    std_logic := 'U';
          BIT_CLK               : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0   : in    std_logic := 'U';
          N_106_mux_i_i         : in    std_logic := 'U';
          TX_collision_detect_i : out   std_logic;
          TX_collision_detect   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component TX_SM
    port( manches_in_dly      : in    std_logic_vector(1 downto 0) := (others => 'U');
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          N_268_i             : out   std_logic;
          N_519               : in    std_logic := 'U';
          N_520               : in    std_logic := 'U';
          N_521               : in    std_logic := 'U';
          N_228               : in    std_logic := 'U';
          N_522               : in    std_logic := 'U';
          N_516               : in    std_logic := 'U';
          N_517               : in    std_logic := 'U';
          N_518               : in    std_logic := 'U';
          TX_FIFO_rd_en       : out   std_logic;
          TX_FIFO_Empty       : in    std_logic := 'U';
          TX_DataEn           : out   std_logic;
          TX_PreAmble         : out   std_logic;
          TX_PostAmble        : out   std_logic;
          tx_crc_byte1_en     : out   std_logic;
          tx_crc_byte2_en     : out   std_logic;
          tx_packet_complt    : out   std_logic;
          iTX_FIFO_rd_en      : out   std_logic;
          start_tx_FIFO       : in    std_logic := 'U';
          DRVR_EN_c           : out   std_logic;
          tx_crc_gen          : out   std_logic;
          byte_clk_en         : in    std_logic := 'U';
          tx_preamble_pat_en  : out   std_logic;
          BIT_CLK             : in    std_logic := 'U';
          N_480_i             : in    std_logic := 'U'
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \MANCH_OUT_P_c\, \byte_clk_en_d[0]_net_1\, VCC_net_1, 
        GND_net_1, \byte_clk_en_d[1]_net_1\, \p2s_data[0]_net_1\, 
        \p2s_data_8[0]\, \p2s_data[1]_net_1\, \p2s_data_8[1]\, 
        \p2s_data[2]_net_1\, \p2s_data_8[2]\, \p2s_data[3]_net_1\, 
        \p2s_data_8[3]\, \p2s_data[4]_net_1\, \p2s_data_8[4]\, 
        \p2s_data[5]_net_1\, \p2s_data_8[5]\, \p2s_data[6]_net_1\, 
        \p2s_data_8[6]\, \p2s_data_0\, \p2s_data_8[7]\, 
        \TX_DataEn_d1\, TX_DataEn, TX_PostAmble, 
        \tx_preamble_pat_en\, p2s_data_8_ss0, tx_crc_byte1_en, 
        \p2s_data_8_m3_0[4]\, \p2s_data_8_m3_0[6]\, 
        \tx_crc_data[8]\, \p2s_data_8_m2_1_1[0]\, 
        \p2s_data_8_m3_0[5]\, \p2s_data_8_m3_0[7]\, 
        \p2s_data_8_m3_0[3]\, \p2s_data_8_m3_0[2]\, 
        \p2s_data_8_m3_0[1]\, \tx_crc_data[14]\, 
        \p2s_data_8_m3_2[6]\, \tx_crc_data[12]\, 
        \p2s_data_8_m3_2[4]\, \tx_crc_data[13]\, 
        \p2s_data_8_m3_2[5]\, \tx_crc_data[10]\, 
        \p2s_data_8_m3_2[2]\, \tx_crc_data[11]\, 
        \p2s_data_8_m3_2[3]\, \tx_crc_data[15]\, 
        \p2s_data_8_m3_2[7]\, \tx_crc_data[9]\, 
        \p2s_data_8_m3_2[1]\, \p2s_data_8_m3_3[7]\, 
        \p2s_data_8_m3_1[7]\, \p2s_data_8_m3_3[4]\, 
        \p2s_data_8_m3_1[4]\, \p2s_data_8_m3_3[3]\, 
        \p2s_data_8_m3_1[3]\, \p2s_data_8_m3_3[2]\, 
        \p2s_data_8_m3_1[2]\, \p2s_data_8_m3_3[1]\, 
        \p2s_data_8_m3_1[1]\, \p2s_data_8_m3_3[5]\, 
        \p2s_data_8_m3_1[5]\, \p2s_data_8_m3_3[6]\, 
        \p2s_data_8_m3_1[6]\, \tx_crc_data[0]\, N_239, 
        \p2s_data_8_m2[0]\, \tx_crc_data[6]\, \tx_crc_data[4]\, 
        \tx_crc_data[5]\, \tx_crc_data[2]\, \tx_crc_data[3]\, 
        \tx_crc_data[7]\, \tx_crc_data[1]\, tx_crc_byte2_en, 
        \DRVR_EN_c\, tx_crc_gen : std_logic;

    for all : CRC16_Generator_0
	Use entity work.CRC16_Generator_0(DEF_ARCH);
    for all : TX_Collision_Detector
	Use entity work.TX_Collision_Detector(DEF_ARCH);
    for all : TX_SM
	Use entity work.TX_SM(DEF_ARCH);
begin 

    p2s_data_0 <= \p2s_data_0\;
    DRVR_EN_c <= \DRVR_EN_c\;
    tx_preamble_pat_en <= \tx_preamble_pat_en\;
    MANCH_OUT_P_c <= \MANCH_OUT_P_c\;

    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_2[4]\ : CFG4
      generic map(INIT => x"3064")

      port map(A => \tx_preamble_pat_en\, B => p2s_data_8_ss0, C
         => \tx_crc_data[12]\, D => tx_crc_byte1_en, Y => 
        \p2s_data_8_m3_2[4]\);
    
    \MAN_OUT_DATA_PROC.un19_tx_dataen\ : CFG2
      generic map(INIT => x"E")

      port map(A => TX_DataEn, B => \TX_DataEn_d1\, Y => 
        un19_tx_dataen);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_3[7]\ : CFG4
      generic map(INIT => x"DDA0")

      port map(A => N_239, B => \tx_crc_data[7]\, C => N_522, D
         => \p2s_data_8_m3_2[7]\, Y => \p2s_data_8_m3_3[7]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_1[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \p2s_data[5]_net_1\, B => N_239, C => 
        \p2s_data_8_m3_0[6]\, Y => \p2s_data_8_m3_1[6]\);
    
    \byte_clk_en_d[0]\ : SLE
      port map(D => byte_clk_en, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => N_480_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \byte_clk_en_d[0]_net_1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8[6]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => TX_DataEn, B => \byte_clk_en_d[0]_net_1\, C
         => \p2s_data_8_m3_3[6]\, D => \p2s_data_8_m3_1[6]\, Y
         => \p2s_data_8[6]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_3[4]\ : CFG4
      generic map(INIT => x"DDA0")

      port map(A => N_239, B => \tx_crc_data[4]\, C => N_520, D
         => \p2s_data_8_m3_2[4]\, Y => \p2s_data_8_m3_3[4]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8[5]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => TX_DataEn, B => \byte_clk_en_d[0]_net_1\, C
         => \p2s_data_8_m3_3[5]\, D => \p2s_data_8_m3_1[5]\, Y
         => \p2s_data_8[5]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8[7]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => TX_DataEn, B => \byte_clk_en_d[0]_net_1\, C
         => \p2s_data_8_m3_3[7]\, D => \p2s_data_8_m3_1[7]\, Y
         => \p2s_data_8[7]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m2[0]\ : CFG4
      generic map(INIT => x"D855")

      port map(A => \p2s_data_8_m2_1_1[0]\, B => N_516, C => 
        \tx_crc_data[0]\, D => N_239, Y => \p2s_data_8_m2[0]\);
    
    \p2s_data[0]\ : SLE
      port map(D => \p2s_data_8[0]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[0]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \p2s_data[6]\ : SLE
      port map(D => \p2s_data_8[6]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[6]_net_1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_0[3]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => \tx_preamble_pat_en\, B => p2s_data_8_ss0, C
         => \p2s_data[2]_net_1\, D => tx_crc_byte1_en, Y => 
        \p2s_data_8_m3_0[3]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_0[7]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => \tx_preamble_pat_en\, B => p2s_data_8_ss0, C
         => \p2s_data[6]_net_1\, D => tx_crc_byte1_en, Y => 
        \p2s_data_8_m3_0[7]\);
    
    \byte_clk_en_d[1]\ : SLE
      port map(D => \byte_clk_en_d[0]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \byte_clk_en_d[1]_net_1\);
    
    TX_CRC_GEN_INST : CRC16_Generator_0
      port map(tx_crc_data(15) => \tx_crc_data[15]\, 
        tx_crc_data(14) => \tx_crc_data[14]\, tx_crc_data(13) => 
        \tx_crc_data[13]\, tx_crc_data(12) => \tx_crc_data[12]\, 
        tx_crc_data(11) => \tx_crc_data[11]\, tx_crc_data(10) => 
        \tx_crc_data[10]\, tx_crc_data(9) => \tx_crc_data[9]\, 
        tx_crc_data(8) => \tx_crc_data[8]\, tx_crc_data(7) => 
        \tx_crc_data[7]\, tx_crc_data(6) => \tx_crc_data[6]\, 
        tx_crc_data(5) => \tx_crc_data[5]\, tx_crc_data(4) => 
        \tx_crc_data[4]\, tx_crc_data(3) => \tx_crc_data[3]\, 
        tx_crc_data(2) => \tx_crc_data[2]\, tx_crc_data(1) => 
        \tx_crc_data[1]\, tx_crc_data(0) => \tx_crc_data[0]\, 
        N_518 => N_518, N_519 => N_519, N_228 => N_228, N_520 => 
        N_520, N_521 => N_521, N_516 => N_516, N_517 => N_517, 
        N_522 => N_522, tx_crc_gen => tx_crc_gen, byte_clk_en => 
        byte_clk_en, BIT_CLK => BIT_CLK, N_9_0_i_i => N_9_0_i_i);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_3[3]\ : CFG4
      generic map(INIT => x"DDA0")

      port map(A => N_239, B => \tx_crc_data[3]\, C => N_519, D
         => \p2s_data_8_m3_2[3]\, Y => \p2s_data_8_m3_3[3]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8[1]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => TX_DataEn, B => \byte_clk_en_d[0]_net_1\, C
         => \p2s_data_8_m3_3[1]\, D => \p2s_data_8_m3_1[1]\, Y
         => \p2s_data_8[1]\);
    
    TX_COLLISION_DETECTOR_INST : TX_Collision_Detector
      port map(p2s_data(7) => \p2s_data_0\, p2s_data(6) => 
        \p2s_data[6]_net_1\, p2s_data(5) => \p2s_data[5]_net_1\, 
        p2s_data(4) => \p2s_data[4]_net_1\, p2s_data(3) => 
        \p2s_data[3]_net_1\, p2s_data(2) => \p2s_data[2]_net_1\, 
        p2s_data(1) => \p2s_data[1]_net_1\, p2s_data(0) => 
        \p2s_data[0]_net_1\, RX_FIFO_DIN(7) => RX_FIFO_DIN(7), 
        RX_FIFO_DIN(6) => RX_FIFO_DIN(6), RX_FIFO_DIN(5) => 
        RX_FIFO_DIN(5), RX_FIFO_DIN(4) => RX_FIFO_DIN(4), 
        RX_FIFO_DIN(3) => RX_FIFO_DIN(3), RX_FIFO_DIN(2) => 
        RX_FIFO_DIN(2), RX_FIFO_DIN(1) => RX_FIFO_DIN(1), 
        RX_FIFO_DIN(0) => RX_FIFO_DIN(0), RX_FIFO_DIN_pipe_0 => 
        RX_FIFO_DIN_pipe_0, byte_clk_en_d_0 => 
        \byte_clk_en_d[1]_net_1\, rx_crc_HighByte_en => 
        rx_crc_HighByte_en, DRVR_EN_c => \DRVR_EN_c\, N_6_0 => 
        N_6_0, tx_col_detect_en => tx_col_detect_en, N_366_i => 
        N_366_i, BIT_CLK => BIT_CLK, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, N_106_mux_i_i => N_106_mux_i_i, 
        TX_collision_detect_i => TX_collision_detect_i, 
        TX_collision_detect => TX_collision_detect);
    
    \p2s_data[2]\ : SLE
      port map(D => \p2s_data_8[2]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[2]_net_1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_0[1]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => \tx_preamble_pat_en\, B => p2s_data_8_ss0, C
         => \p2s_data[0]_net_1\, D => tx_crc_byte1_en, Y => 
        \p2s_data_8_m3_0[1]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_3[6]\ : CFG4
      generic map(INIT => x"DDA0")

      port map(A => N_239, B => \tx_crc_data[6]\, C => N_228, D
         => \p2s_data_8_m3_2[6]\, Y => \p2s_data_8_m3_3[6]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_2[5]\ : CFG4
      generic map(INIT => x"3064")

      port map(A => \tx_preamble_pat_en\, B => p2s_data_8_ss0, C
         => \tx_crc_data[13]\, D => tx_crc_byte1_en, Y => 
        \p2s_data_8_m3_2[5]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \TX_PostAmble_d1\ : SLE
      port map(D => TX_PostAmble, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => N_480_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => TX_PostAmble_d1);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_2[3]\ : CFG4
      generic map(INIT => x"3064")

      port map(A => \tx_preamble_pat_en\, B => p2s_data_8_ss0, C
         => \tx_crc_data[11]\, D => tx_crc_byte1_en, Y => 
        \p2s_data_8_m3_2[3]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_0[5]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => \tx_preamble_pat_en\, B => p2s_data_8_ss0, C
         => \p2s_data[4]_net_1\, D => tx_crc_byte1_en, Y => 
        \p2s_data_8_m3_0[5]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_0[2]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => \tx_preamble_pat_en\, B => p2s_data_8_ss0, C
         => \p2s_data[1]_net_1\, D => tx_crc_byte1_en, Y => 
        \p2s_data_8_m3_0[2]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_1[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \p2s_data[0]_net_1\, B => N_239, C => 
        \p2s_data_8_m3_0[1]\, Y => \p2s_data_8_m3_1[1]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8[2]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => TX_DataEn, B => \byte_clk_en_d[0]_net_1\, C
         => \p2s_data_8_m3_3[2]\, D => \p2s_data_8_m3_1[2]\, Y
         => \p2s_data_8[2]\);
    
    \p2s_data[4]\ : SLE
      port map(D => \p2s_data_8[4]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[4]_net_1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_2[1]\ : CFG4
      generic map(INIT => x"3064")

      port map(A => \tx_preamble_pat_en\, B => p2s_data_8_ss0, C
         => \tx_crc_data[9]\, D => tx_crc_byte1_en, Y => 
        \p2s_data_8_m3_2[1]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_1[5]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \p2s_data[4]_net_1\, B => N_239, C => 
        \p2s_data_8_m3_0[5]\, Y => \p2s_data_8_m3_1[5]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_1[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \p2s_data[3]_net_1\, B => N_239, C => 
        \p2s_data_8_m3_0[4]\, Y => \p2s_data_8_m3_1[4]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_2[2]\ : CFG4
      generic map(INIT => x"3064")

      port map(A => \tx_preamble_pat_en\, B => p2s_data_8_ss0, C
         => \tx_crc_data[10]\, D => tx_crc_byte1_en, Y => 
        \p2s_data_8_m3_2[2]\);
    
    TRANSMIT_SM : TX_SM
      port map(manches_in_dly(1) => manches_in_dly(1), 
        manches_in_dly(0) => manches_in_dly(0), 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, N_268_i => 
        N_268_i, N_519 => N_519, N_520 => N_520, N_521 => N_521, 
        N_228 => N_228, N_522 => N_522, N_516 => N_516, N_517 => 
        N_517, N_518 => N_518, TX_FIFO_rd_en => TX_FIFO_rd_en, 
        TX_FIFO_Empty => TX_FIFO_Empty, TX_DataEn => TX_DataEn, 
        TX_PreAmble => TX_PreAmble, TX_PostAmble => TX_PostAmble, 
        tx_crc_byte1_en => tx_crc_byte1_en, tx_crc_byte2_en => 
        tx_crc_byte2_en, tx_packet_complt => tx_packet_complt, 
        iTX_FIFO_rd_en => iTX_FIFO_rd_en, start_tx_FIFO => 
        start_tx_FIFO, DRVR_EN_c => \DRVR_EN_c\, tx_crc_gen => 
        tx_crc_gen, byte_clk_en => byte_clk_en, 
        tx_preamble_pat_en => \tx_preamble_pat_en\, BIT_CLK => 
        BIT_CLK, N_480_i => N_480_i);
    
    \p2s_data[1]\ : SLE
      port map(D => \p2s_data_8[1]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[1]_net_1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_3[5]\ : CFG4
      generic map(INIT => x"DDA0")

      port map(A => N_239, B => \tx_crc_data[5]\, C => N_521, D
         => \p2s_data_8_m3_2[5]\, Y => \p2s_data_8_m3_3[5]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_1[2]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \p2s_data[1]_net_1\, B => N_239, C => 
        \p2s_data_8_m3_0[2]\, Y => \p2s_data_8_m3_1[2]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_0[6]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => \tx_preamble_pat_en\, B => p2s_data_8_ss0, C
         => \p2s_data[5]_net_1\, D => tx_crc_byte1_en, Y => 
        \p2s_data_8_m3_0[6]\);
    
    \p2s_data[3]\ : SLE
      port map(D => \p2s_data_8[3]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[3]_net_1\);
    
    MANCHESTER_OUT : SLE
      port map(D => MANCHESTER_OUT_5, CLK => CommsFPGA_CCC_0_GL1, 
        EN => VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \MANCH_OUT_P_c\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m2_1_1[0]\ : CFG4
      generic map(INIT => x"0313")

      port map(A => \tx_preamble_pat_en\, B => p2s_data_8_ss0, C
         => \tx_crc_data[8]\, D => tx_crc_byte1_en, Y => 
        \p2s_data_8_m2_1_1[0]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m2s2_i_a5\ : CFG2
      generic map(INIT => x"1")

      port map(A => \tx_preamble_pat_en\, B => tx_crc_byte1_en, Y
         => N_239);
    
    MANCHESTER_OUT_RNI19ND : CFG1
      generic map(INIT => "01")

      port map(A => \MANCH_OUT_P_c\, Y => MANCH_OUT_P_c_i);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_3[1]\ : CFG4
      generic map(INIT => x"DDA0")

      port map(A => N_239, B => \tx_crc_data[1]\, C => N_517, D
         => \p2s_data_8_m3_2[1]\, Y => \p2s_data_8_m3_3[1]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_3[2]\ : CFG4
      generic map(INIT => x"DDA0")

      port map(A => N_239, B => \tx_crc_data[2]\, C => N_518, D
         => \p2s_data_8_m3_2[2]\, Y => \p2s_data_8_m3_3[2]\);
    
    \p2s_data[5]\ : SLE
      port map(D => \p2s_data_8[5]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[5]_net_1\);
    
    TX_DataEn_d1 : SLE
      port map(D => TX_DataEn, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => N_480_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \TX_DataEn_d1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_1[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \p2s_data[6]_net_1\, B => N_239, C => 
        \p2s_data_8_m3_0[7]\, Y => \p2s_data_8_m3_1[7]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8[0]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \byte_clk_en_d[0]_net_1\, B => TX_DataEn, C
         => \p2s_data_8_m2[0]\, Y => \p2s_data_8[0]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8[4]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => TX_DataEn, B => \byte_clk_en_d[0]_net_1\, C
         => \p2s_data_8_m3_3[4]\, D => \p2s_data_8_m3_1[4]\, Y
         => \p2s_data_8[4]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_0[4]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => \tx_preamble_pat_en\, B => p2s_data_8_ss0, C
         => \p2s_data[3]_net_1\, D => tx_crc_byte1_en, Y => 
        \p2s_data_8_m3_0[4]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8[3]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => TX_DataEn, B => \byte_clk_en_d[0]_net_1\, C
         => \p2s_data_8_m3_3[3]\, D => \p2s_data_8_m3_1[3]\, Y
         => \p2s_data_8[3]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_2[6]\ : CFG4
      generic map(INIT => x"3064")

      port map(A => \tx_preamble_pat_en\, B => p2s_data_8_ss0, C
         => \tx_crc_data[14]\, D => tx_crc_byte1_en, Y => 
        \p2s_data_8_m3_2[6]\);
    
    \p2s_data[7]\ : SLE
      port map(D => \p2s_data_8[7]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data_0\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_ss0_0_o5\ : CFG3
      generic map(INIT => x"DC")

      port map(A => tx_crc_byte1_en, B => \tx_preamble_pat_en\, C
         => tx_crc_byte2_en, Y => p2s_data_8_ss0);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_2[7]\ : CFG4
      generic map(INIT => x"FCEC")

      port map(A => \tx_preamble_pat_en\, B => p2s_data_8_ss0, C
         => \tx_crc_data[15]\, D => tx_crc_byte1_en, Y => 
        \p2s_data_8_m3_2[7]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_8_m3_1[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \p2s_data[2]_net_1\, B => N_239, C => 
        \p2s_data_8_m3_0[3]\, Y => \p2s_data_8_m3_1[3]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity IdleLineDetectorZ1 is

    port( N_268_i             : in    std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          N_480_i             : in    std_logic;
          idle_line           : out   std_logic
        );

end IdleLineDetectorZ1;

architecture DEF_ARCH of IdleLineDetectorZ1 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, N_341_i, GND_net_1, 
        \idle_line_cntr[0]_net_1\, \idle_line_cntr_s[0]\, 
        \idle_line_cntr[1]_net_1\, \idle_line_cntr_s[1]\, 
        \idle_line_cntr[2]_net_1\, \idle_line_cntr_s[2]\, 
        \idle_line_cntr[3]_net_1\, \idle_line_cntr_s[3]\, 
        \idle_line_cntr[4]_net_1\, \idle_line_cntr_s[4]\, 
        \idle_line_cntr[5]_net_1\, \idle_line_cntr_s[5]_net_1\, 
        idle_line_cntr_cry_cy, \idle_line_cntr_cry_cy_Y_0[0]\, 
        un5_manches_in_dly_3, \idle_line_cntr_cry[0]_net_1\, 
        \idle_line_cntr_cry[1]_net_1\, 
        \idle_line_cntr_cry[2]_net_1\, 
        \idle_line_cntr_cry[3]_net_1\, 
        \idle_line_cntr_cry[4]_net_1\ : std_logic;

begin 


    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_3_RNI1QPI\ : CFG4
      generic map(INIT => x"2000")

      port map(A => un5_manches_in_dly_3, B => N_268_i, C => 
        \idle_line_cntr[5]_net_1\, D => \idle_line_cntr[4]_net_1\, 
        Y => N_341_i);
    
    \idle_line_cntr_cry[2]\ : ARI1
      generic map(INIT => x"4AC00")

      port map(A => VCC_net_1, B => \idle_line_cntr[2]_net_1\, C
         => N_341_i, D => \idle_line_cntr_cry_cy_Y_0[0]\, FCI => 
        \idle_line_cntr_cry[1]_net_1\, S => \idle_line_cntr_s[2]\, 
        Y => OPEN, FCO => \idle_line_cntr_cry[2]_net_1\);
    
    \idle_line_cntr_s[5]\ : ARI1
      generic map(INIT => x"4AC00")

      port map(A => VCC_net_1, B => \idle_line_cntr[5]_net_1\, C
         => N_341_i, D => \idle_line_cntr_cry_cy_Y_0[0]\, FCI => 
        \idle_line_cntr_cry[4]_net_1\, S => 
        \idle_line_cntr_s[5]_net_1\, Y => OPEN, FCO => OPEN);
    
    \idle_line_cntr[0]\ : SLE
      port map(D => \idle_line_cntr_s[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[0]_net_1\);
    
    \idle_line\ : SLE
      port map(D => N_341_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        idle_line);
    
    \idle_line_cntr_cry[4]\ : ARI1
      generic map(INIT => x"4AC00")

      port map(A => VCC_net_1, B => \idle_line_cntr[4]_net_1\, C
         => N_341_i, D => \idle_line_cntr_cry_cy_Y_0[0]\, FCI => 
        \idle_line_cntr_cry[3]_net_1\, S => \idle_line_cntr_s[4]\, 
        Y => OPEN, FCO => \idle_line_cntr_cry[4]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \idle_line_cntr_cry[0]\ : ARI1
      generic map(INIT => x"4AC00")

      port map(A => VCC_net_1, B => \idle_line_cntr[0]_net_1\, C
         => N_341_i, D => \idle_line_cntr_cry_cy_Y_0[0]\, FCI => 
        idle_line_cntr_cry_cy, S => \idle_line_cntr_s[0]\, Y => 
        OPEN, FCO => \idle_line_cntr_cry[0]_net_1\);
    
    \idle_line_cntr_cry[3]\ : ARI1
      generic map(INIT => x"4AC00")

      port map(A => VCC_net_1, B => \idle_line_cntr[3]_net_1\, C
         => N_341_i, D => \idle_line_cntr_cry_cy_Y_0[0]\, FCI => 
        \idle_line_cntr_cry[2]_net_1\, S => \idle_line_cntr_s[3]\, 
        Y => OPEN, FCO => \idle_line_cntr_cry[3]_net_1\);
    
    \idle_line_cntr_cry_cy[0]\ : ARI1
      generic map(INIT => x"4007F")

      port map(A => N_268_i, B => un5_manches_in_dly_3, C => 
        \idle_line_cntr[4]_net_1\, D => \idle_line_cntr[5]_net_1\, 
        FCI => VCC_net_1, S => OPEN, Y => 
        \idle_line_cntr_cry_cy_Y_0[0]\, FCO => 
        idle_line_cntr_cry_cy);
    
    \idle_line_cntr_cry[1]\ : ARI1
      generic map(INIT => x"4AC00")

      port map(A => VCC_net_1, B => \idle_line_cntr[1]_net_1\, C
         => N_341_i, D => \idle_line_cntr_cry_cy_Y_0[0]\, FCI => 
        \idle_line_cntr_cry[0]_net_1\, S => \idle_line_cntr_s[1]\, 
        Y => OPEN, FCO => \idle_line_cntr_cry[1]_net_1\);
    
    \idle_line_cntr[4]\ : SLE
      port map(D => \idle_line_cntr_s[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[4]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \idle_line_cntr[5]\ : SLE
      port map(D => \idle_line_cntr_s[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[5]_net_1\);
    
    \idle_line_cntr[1]\ : SLE
      port map(D => \idle_line_cntr_s[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[1]_net_1\);
    
    \idle_line_cntr[3]\ : SLE
      port map(D => \idle_line_cntr_s[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[3]_net_1\);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_3\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \idle_line_cntr[3]_net_1\, B => 
        \idle_line_cntr[2]_net_1\, C => \idle_line_cntr[1]_net_1\, 
        D => \idle_line_cntr[0]_net_1\, Y => un5_manches_in_dly_3);
    
    \idle_line_cntr[2]\ : SLE
      port map(D => \idle_line_cntr_s[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[2]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity ManchesDecoder_Adapter is

    port( manches_in_dly      : out   std_logic_vector(1 downto 0);
          RX_FIFO_DIN         : out   std_logic_vector(7 downto 0);
          idle_line           : out   std_logic;
          N_268_i             : in    std_logic;
          internal_loopback   : in    std_logic;
          MANCHESTER_IN_c     : in    std_logic;
          MANCH_OUT_P_c       : in    std_logic;
          irx_center_sample   : out   std_logic;
          N_447_i_i           : in    std_logic;
          sampler_clk1x_en    : out   std_logic;
          N_480_i             : in    std_logic;
          clk1x_enable        : in    std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          N_584_i_i           : in    std_logic
        );

end ManchesDecoder_Adapter;

architecture DEF_ARCH of ManchesDecoder_Adapter is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IdleLineDetectorZ1
    port( N_268_i             : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          N_480_i             : in    std_logic := 'U';
          idle_line           : out   std_logic
        );
  end component;

    signal \clock_adjust\, clock_adjust_i, \clkdiv[2]_net_1\, 
        VCC_net_1, N_327_i_i, GND_net_1, \clkdiv[3]_net_1\, 
        N_352_i_i, \decoder_Transition_d[0]_net_1\, 
        \decoder_Transition\, \decoder_Transition_d[1]_net_1\, 
        \decoder_Transition_d[2]_net_1\, \RX_FIFO_DIN[0]\, 
        \iNRZ_data\, \sampler_clk1x_en\, \RX_FIFO_DIN[1]\, 
        \RX_FIFO_DIN[2]\, \RX_FIFO_DIN[3]\, \RX_FIFO_DIN[4]\, 
        \RX_FIFO_DIN[5]\, \RX_FIFO_DIN[6]\, \manches_in_dly[0]\, 
        \un1_manches_in[0]_net_1\, \manches_in_dly[1]\, 
        \clkdiv[0]_net_1\, N_306_i, \clkdiv[1]_net_1\, N_315_i_i, 
        \decoder_ShiftReg[0]_net_1\, \manches_ShiftReg[0]_net_1\, 
        N_305_i, irx_center_sample_net_1, isampler_clk1x_en_1, 
        decoder_Transition_1, \manches_Transition\, 
        manches_Transition_1, un16_irx_center_sample, 
        un16_clk1x_enable, N_274 : std_logic;

    for all : IdleLineDetectorZ1
	Use entity work.IdleLineDetectorZ1(DEF_ARCH);
begin 

    manches_in_dly(1) <= \manches_in_dly[1]\;
    manches_in_dly(0) <= \manches_in_dly[0]\;
    RX_FIFO_DIN(6) <= \RX_FIFO_DIN[6]\;
    RX_FIFO_DIN(5) <= \RX_FIFO_DIN[5]\;
    RX_FIFO_DIN(4) <= \RX_FIFO_DIN[4]\;
    RX_FIFO_DIN(3) <= \RX_FIFO_DIN[3]\;
    RX_FIFO_DIN(2) <= \RX_FIFO_DIN[2]\;
    RX_FIFO_DIN(1) <= \RX_FIFO_DIN[1]\;
    RX_FIFO_DIN(0) <= \RX_FIFO_DIN[0]\;
    irx_center_sample <= irx_center_sample_net_1;
    sampler_clk1x_en <= \sampler_clk1x_en\;

    \un1_clkdiv_1.SUM_0_x2[0]\ : CFG3
      generic map(INIT => x"A6")

      port map(A => \clkdiv[0]_net_1\, B => clk1x_enable, C => 
        \clock_adjust\, Y => N_306_i);
    
    \s2p_data[2]\ : SLE
      port map(D => \RX_FIFO_DIN[1]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => N_480_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[2]\);
    
    \imanches_in_dly[0]\ : SLE
      port map(D => \un1_manches_in[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \manches_in_dly[0]\);
    
    \un1_clkdiv_1.SUM_0_o2[1]\ : CFG3
      generic map(INIT => x"F7")

      port map(A => \clkdiv[0]_net_1\, B => clk1x_enable, C => 
        \clock_adjust\, Y => N_274);
    
    \decoder_Transition_d[2]\ : SLE
      port map(D => \decoder_Transition_d[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => N_584_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \decoder_Transition_d[2]_net_1\);
    
    \NRZ_DATA_PROC.iNRZ_data_1_0_x2\ : CFG2
      generic map(INIT => x"6")

      port map(A => \manches_in_dly[1]\, B => \clkdiv[3]_net_1\, 
        Y => N_305_i);
    
    \un1_clkdiv_1.N_327_i_i\ : CFG3
      generic map(INIT => x"D2")

      port map(A => \clkdiv[1]_net_1\, B => N_274, C => 
        \clkdiv[2]_net_1\, Y => N_327_i_i);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \s2p_data[4]\ : SLE
      port map(D => \RX_FIFO_DIN[3]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => N_480_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[4]\);
    
    clock_adjust_RNIMA1A : CFG1
      generic map(INIT => "01")

      port map(A => \clock_adjust\, Y => clock_adjust_i);
    
    \irx_center_sample\ : SLE
      port map(D => un16_irx_center_sample, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clock_adjust_i, ALn => N_480_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => irx_center_sample_net_1);
    
    \s2p_data[1]\ : SLE
      port map(D => \RX_FIFO_DIN[0]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => N_480_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[1]\);
    
    \decoder_ShiftReg[0]\ : SLE
      port map(D => \clkdiv[3]_net_1\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => clk1x_enable, ALn => N_584_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \decoder_ShiftReg[0]_net_1\);
    
    \manches_ShiftReg[0]\ : SLE
      port map(D => \manches_in_dly[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => N_584_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \manches_ShiftReg[0]_net_1\);
    
    iNRZ_data : SLE
      port map(D => N_305_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        irx_center_sample_net_1, ALn => N_447_i_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \iNRZ_data\);
    
    \clkdiv[2]\ : SLE
      port map(D => N_327_i_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => N_584_i_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \clkdiv[2]_net_1\);
    
    \s2p_data[3]\ : SLE
      port map(D => \RX_FIFO_DIN[2]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => N_480_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[3]\);
    
    \decoder_Transition_d[0]\ : SLE
      port map(D => \decoder_Transition\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => N_584_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \decoder_Transition_d[0]_net_1\);
    
    decoder_Transition : SLE
      port map(D => decoder_Transition_1, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => N_584_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \decoder_Transition\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \clkdiv[1]\ : SLE
      port map(D => N_315_i_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => N_584_i_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \clkdiv[1]_net_1\);
    
    \s2p_data[5]\ : SLE
      port map(D => \RX_FIFO_DIN[4]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => N_480_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[5]\);
    
    \un1_clkdiv_1.N_315_i_i\ : CFG4
      generic map(INIT => x"B4F0")

      port map(A => \clock_adjust\, B => \clkdiv[0]_net_1\, C => 
        \clkdiv[1]_net_1\, D => clk1x_enable, Y => N_315_i_i);
    
    RX_IDLE_LINE_DETECTOR : IdleLineDetectorZ1
      port map(N_268_i => N_268_i, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, N_480_i => N_480_i, idle_line => 
        idle_line);
    
    un10_clk1x_enable : CFG2
      generic map(INIT => x"6")

      port map(A => \clkdiv[3]_net_1\, B => 
        \decoder_ShiftReg[0]_net_1\, Y => decoder_Transition_1);
    
    \RX_CENTER_SAMPLE_PROC.un16_irx_center_sample_0_a2\ : CFG3
      generic map(INIT => x"40")

      port map(A => \clkdiv[2]_net_1\, B => \clkdiv[1]_net_1\, C
         => \clkdiv[0]_net_1\, Y => un16_irx_center_sample);
    
    clock_adjust : SLE
      port map(D => un16_clk1x_enable, CLK => CommsFPGA_CCC_0_GL0, 
        EN => clk1x_enable, ALn => N_584_i_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \clock_adjust\);
    
    \un1_manches_in[0]\ : CFG3
      generic map(INIT => x"A3")

      port map(A => MANCH_OUT_P_c, B => MANCHESTER_IN_c, C => 
        internal_loopback, Y => \un1_manches_in[0]_net_1\);
    
    \SAMPLE_CLK1X_EN_PROC.isampler_clk1x_en_1_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \clkdiv[0]_net_1\, B => \clkdiv[3]_net_1\, C
         => \clkdiv[2]_net_1\, D => \clkdiv[1]_net_1\, Y => 
        isampler_clk1x_en_1);
    
    manches_Transition : SLE
      port map(D => manches_Transition_1, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => N_584_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \manches_Transition\);
    
    \un1_clkdiv_1.N_352_i_i\ : CFG4
      generic map(INIT => x"F708")

      port map(A => \clkdiv[1]_net_1\, B => \clkdiv[2]_net_1\, C
         => N_274, D => \clkdiv[3]_net_1\, Y => N_352_i_i);
    
    \CLOCK_ADJUST_PROC.un16_clk1x_enable\ : CFG2
      generic map(INIT => x"8")

      port map(A => \decoder_Transition_d[2]_net_1\, B => 
        \manches_Transition\, Y => un16_clk1x_enable);
    
    \s2p_data[7]\ : SLE
      port map(D => \RX_FIFO_DIN[6]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => N_480_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RX_FIFO_DIN(7));
    
    \clkdiv[0]\ : SLE
      port map(D => N_306_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => N_584_i_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \clkdiv[0]_net_1\);
    
    \clkdiv[3]\ : SLE
      port map(D => N_352_i_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => N_584_i_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \clkdiv[3]_net_1\);
    
    \imanches_in_dly[1]\ : SLE
      port map(D => \manches_in_dly[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \manches_in_dly[1]\);
    
    \decoder_Transition_d[1]\ : SLE
      port map(D => \decoder_Transition_d[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => N_584_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \decoder_Transition_d[1]_net_1\);
    
    \s2p_data[0]\ : SLE
      port map(D => \iNRZ_data\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \sampler_clk1x_en\, ALn => N_480_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RX_FIFO_DIN[0]\);
    
    \s2p_data[6]\ : SLE
      port map(D => \RX_FIFO_DIN[5]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => N_480_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[6]\);
    
    un4_clk1x_enable : CFG2
      generic map(INIT => x"6")

      port map(A => \manches_in_dly[1]\, B => 
        \manches_ShiftReg[0]_net_1\, Y => manches_Transition_1);
    
    isampler_clk1x_en : SLE
      port map(D => isampler_clk1x_en_1, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clock_adjust_i, ALn => N_480_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \sampler_clk1x_en\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CRC16_Generator_1 is

    port( RX_FIFO_DIN         : in    std_logic_vector(7 downto 0);
          rx_crc_data_calc    : out   std_logic_vector(15 downto 0);
          rx_crc_gen          : in    std_logic;
          sampler_clk1x_en    : in    std_logic;
          iRX_FIFO_wr_en      : in    std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          rx_crc_reset_i      : in    std_logic
        );

end CRC16_Generator_1;

architecture DEF_ARCH of CRC16_Generator_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \rx_crc_data_calc[13]\, GND_net_1, 
        \rx_crc_data_calc[5]\, \N_343_i\, VCC_net_1, 
        \rx_crc_data_calc[14]\, \rx_crc_data_calc[6]\, 
        \rx_crc_data_calc[15]\, \lfsr_c[15]\, 
        \rx_crc_data_calc[0]\, \lfsr_c[0]\, \rx_crc_data_calc[1]\, 
        \lfsr_c[1]\, \rx_crc_data_calc[2]\, N_316_i, 
        \rx_crc_data_calc[3]\, N_323_i, \rx_crc_data_calc[4]\, 
        N_320_i, N_319_i, N_317_i, \rx_crc_data_calc[7]\, N_318_i, 
        \rx_crc_data_calc[8]\, N_329_i_i, \rx_crc_data_calc[9]\, 
        N_324_i_i, \rx_crc_data_calc[10]\, \rx_crc_data_calc[11]\, 
        \rx_crc_data_calc[12]\, N_263_i : std_logic;

begin 

    rx_crc_data_calc(15) <= \rx_crc_data_calc[15]\;
    rx_crc_data_calc(14) <= \rx_crc_data_calc[14]\;
    rx_crc_data_calc(13) <= \rx_crc_data_calc[13]\;
    rx_crc_data_calc(12) <= \rx_crc_data_calc[12]\;
    rx_crc_data_calc(11) <= \rx_crc_data_calc[11]\;
    rx_crc_data_calc(10) <= \rx_crc_data_calc[10]\;
    rx_crc_data_calc(9) <= \rx_crc_data_calc[9]\;
    rx_crc_data_calc(8) <= \rx_crc_data_calc[8]\;
    rx_crc_data_calc(7) <= \rx_crc_data_calc[7]\;
    rx_crc_data_calc(6) <= \rx_crc_data_calc[6]\;
    rx_crc_data_calc(5) <= \rx_crc_data_calc[5]\;
    rx_crc_data_calc(4) <= \rx_crc_data_calc[4]\;
    rx_crc_data_calc(3) <= \rx_crc_data_calc[3]\;
    rx_crc_data_calc(2) <= \rx_crc_data_calc[2]\;
    rx_crc_data_calc(1) <= \rx_crc_data_calc[1]\;
    rx_crc_data_calc(0) <= \rx_crc_data_calc[0]\;

    \lfsr_q[9]\ : SLE
      port map(D => N_324_i_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_343_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[9]\);
    
    \lfsr_c_0_a2_2_x2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[9]\, B => 
        \rx_crc_data_calc[8]\, C => RX_FIFO_DIN(1), D => 
        RX_FIFO_DIN(0), Y => N_316_i);
    
    N_343_i : CFG3
      generic map(INIT => x"80")

      port map(A => iRX_FIFO_wr_en, B => sampler_clk1x_en, C => 
        rx_crc_gen, Y => \N_343_i\);
    
    \lfsr_q[6]\ : SLE
      port map(D => N_317_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_343_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[6]\);
    
    \lfsr_q[3]\ : SLE
      port map(D => N_323_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_343_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[3]\);
    
    \lfsr_c_0_a2_2_x2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[13]\, B => 
        \rx_crc_data_calc[12]\, C => RX_FIFO_DIN(5), D => 
        RX_FIFO_DIN(4), Y => N_317_i);
    
    \lfsr_q[10]\ : SLE
      port map(D => \rx_crc_data_calc[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \N_343_i\, ALn => 
        rx_crc_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[10]\);
    
    \lfsr_q[2]\ : SLE
      port map(D => N_316_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_343_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[2]\);
    
    \lfsr_c_0_a2_0_x2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[13]\, B => 
        \rx_crc_data_calc[14]\, C => RX_FIFO_DIN(6), D => 
        RX_FIFO_DIN(5), Y => N_318_i);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \lfsr_q[1]\ : SLE
      port map(D => \lfsr_c[1]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \N_343_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rx_crc_data_calc[1]\);
    
    \lfsr_q[7]\ : SLE
      port map(D => N_318_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_343_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[7]\);
    
    \lfsr_c_0_a2_0_x2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[10]\, B => 
        \rx_crc_data_calc[9]\, C => RX_FIFO_DIN(2), D => 
        RX_FIFO_DIN(1), Y => N_323_i);
    
    \lfsr_q[4]\ : SLE
      port map(D => N_320_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_343_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[4]\);
    
    \lfsr_q[11]\ : SLE
      port map(D => \rx_crc_data_calc[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \N_343_i\, ALn => 
        rx_crc_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[11]\);
    
    \lfsr_q[5]\ : SLE
      port map(D => N_319_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_343_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[5]\);
    
    \lfsr_c_0_a2[1]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => N_263_i, B => N_319_i, C => N_318_i, D => 
        N_323_i, Y => \lfsr_c[1]\);
    
    \lfsr_q_RNO[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => N_263_i, B => \rx_crc_data_calc[1]\, Y => 
        N_324_i_i);
    
    \lfsr_q[0]\ : SLE
      port map(D => \lfsr_c[0]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \N_343_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rx_crc_data_calc[0]\);
    
    \lfsr_c_0_a2[15]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[7]\, B => 
        \rx_crc_data_calc[8]\, C => RX_FIFO_DIN(0), D => 
        \lfsr_c[1]\, Y => \lfsr_c[15]\);
    
    \lfsr_q[12]\ : SLE
      port map(D => \rx_crc_data_calc[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \N_343_i\, ALn => 
        rx_crc_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[12]\);
    
    \lfsr_q[14]\ : SLE
      port map(D => \rx_crc_data_calc[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \N_343_i\, ALn => 
        rx_crc_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[14]\);
    
    \lfsr_c_0_a2_i_x2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[14]\, B => 
        \rx_crc_data_calc[0]\, C => N_263_i, D => RX_FIFO_DIN(6), 
        Y => N_329_i_i);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \lfsr_c_0_a2_0_x2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[12]\, B => 
        \rx_crc_data_calc[11]\, C => RX_FIFO_DIN(4), D => 
        RX_FIFO_DIN(3), Y => N_319_i);
    
    \lfsr_c_0_a2_2_x2[4]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[11]\, B => 
        \rx_crc_data_calc[10]\, C => RX_FIFO_DIN(3), D => 
        RX_FIFO_DIN(2), Y => N_320_i);
    
    \lfsr_c_0_a2_1_0_x2[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => RX_FIFO_DIN(7), B => \rx_crc_data_calc[15]\, 
        Y => N_263_i);
    
    \lfsr_q[8]\ : SLE
      port map(D => N_329_i_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_343_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[8]\);
    
    \lfsr_q[13]\ : SLE
      port map(D => \rx_crc_data_calc[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \N_343_i\, ALn => 
        rx_crc_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[13]\);
    
    \lfsr_c_0_a2[0]\ : CFG3
      generic map(INIT => x"96")

      port map(A => RX_FIFO_DIN(0), B => \lfsr_c[1]\, C => 
        \rx_crc_data_calc[8]\, Y => \lfsr_c[0]\);
    
    \lfsr_q[15]\ : SLE
      port map(D => \lfsr_c[15]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \N_343_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rx_crc_data_calc[15]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity ReadFIFO_Write_SM is

    port( consumer_type4_reg                 : in    std_logic_vector(9 downto 0);
          consumer_type3_reg                 : in    std_logic_vector(9 downto 0);
          consumer_type2_reg                 : in    std_logic_vector(9 downto 0);
          consumer_type1_reg                 : in    std_logic_vector(9 downto 0);
          RX_FIFO_DIN                        : in    std_logic_vector(7 downto 0);
          RX_FIFO_DIN_pipe                   : out   std_logic_vector(8 downto 0);
          DRVR_EN_c                          : in    std_logic;
          N_366_i                            : out   std_logic;
          clk1x_enable                       : in    std_logic;
          N_480                              : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY_i_m_i : out   std_logic;
          CoreAPB3_0_APBmslave0_PREADY       : in    std_logic;
          CoreAPB3_0_APBmslave0_PSELx        : in    std_logic;
          tx_col_detect_en                   : in    std_logic;
          TX_collision_detect                : in    std_logic;
          sampler_clk1x_en                   : in    std_logic;
          idle_line                          : in    std_logic;
          packet_avail                       : in    std_logic;
          N_447_i_i                          : out   std_logic;
          RX_InProcess_d1                    : out   std_logic;
          iRX_FIFO_wr_en                     : out   std_logic;
          RX_EarlyTerm                       : out   std_logic;
          rx_crc_HighByte_en                 : out   std_logic;
          CommsFPGA_CCC_0_GL0                : in    std_logic;
          N_480_i                            : in    std_logic;
          rx_packet_complt_i                 : out   std_logic;
          rx_packet_complt                   : out   std_logic;
          rx_CRC_error_i                     : out   std_logic;
          rx_CRC_error                       : out   std_logic
        );

end ReadFIFO_Write_SM;

architecture DEF_ARCH of ReadFIFO_Write_SM is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CRC16_Generator_1
    port( RX_FIFO_DIN         : in    std_logic_vector(7 downto 0) := (others => 'U');
          rx_crc_data_calc    : out   std_logic_vector(15 downto 0);
          rx_crc_gen          : in    std_logic := 'U';
          sampler_clk1x_en    : in    std_logic := 'U';
          iRX_FIFO_wr_en      : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          rx_crc_reset_i      : in    std_logic := 'U'
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal rx_crc_reset_i, \rx_crc_reset\, un8_rst, un8_rst_i, 
        rx_CRC_error_net_1, rx_packet_complt_net_1, 
        \consumer_type[8]_net_1\, VCC_net_1, 
        \consumer_type_12[8]\, N_333_i, GND_net_1, 
        \consumer_type[9]_net_1\, \consumer_type_12[9]\, 
        \SM_advancebit_cntr[0]_net_1\, N_321_i_i, 
        \SM_advancebit_cntr[1]_net_1\, N_325_i_i, 
        \SM_advancebit_cntr[2]_net_1\, N_348_i_i, 
        \bit_cntr[0]_net_1\, un15_rst_i, N_322_i_i, 
        \bit_cntr[1]_net_1\, N_326_i_i, \bit_cntr[2]_net_1\, 
        N_350_i_i, \rx_crc_data_store[9]_net_1\, 
        \RX_FIFO_DIN_pipe[1]\, N_344_i, 
        \rx_crc_data_store[10]_net_1\, \RX_FIFO_DIN_pipe[2]\, 
        \rx_crc_data_store[11]_net_1\, \RX_FIFO_DIN_pipe[3]\, 
        \rx_crc_data_store[12]_net_1\, \RX_FIFO_DIN_pipe[4]\, 
        \rx_crc_data_store[13]_net_1\, \RX_FIFO_DIN_pipe[5]\, 
        \rx_crc_data_store[14]_net_1\, \RX_FIFO_DIN_pipe[6]\, 
        \rx_crc_data_store[15]_net_1\, \RX_FIFO_DIN_pipe[7]\, 
        \consumer_type[0]_net_1\, \consumer_type_12[0]\, 
        \consumer_type[1]_net_1\, \consumer_type_12[1]\, 
        \consumer_type[2]_net_1\, \consumer_type_12[2]\, 
        \consumer_type[3]_net_1\, \consumer_type_12[3]\, 
        \consumer_type[4]_net_1\, \consumer_type_12[4]\, 
        \consumer_type[5]_net_1\, \consumer_type_12[5]\, 
        \consumer_type[6]_net_1\, \consumer_type_12[6]\, 
        \consumer_type[7]_net_1\, \consumer_type_12[7]\, 
        \rx_packet_length[5]_net_1\, 
        \rx_packet_length_13[5]_net_1\, 
        \un1_ReadFIFO_WR_STATE_14_0_0\, 
        \rx_packet_length[6]_net_1\, 
        \rx_packet_length_13[6]_net_1\, 
        \rx_packet_length[7]_net_1\, 
        \rx_packet_length_13[7]_net_1\, 
        \rx_packet_length[8]_net_1\, N_337_i, 
        \rx_packet_length[9]_net_1\, N_123_i, 
        \rx_packet_length[10]_net_1\, N_125_i, 
        \rx_crc_data_store[0]_net_1\, 
        \un1_rx_fifo_din_d3[0]_net_1\, N_330_i, 
        \rx_crc_data_store[1]_net_1\, 
        \un1_rx_fifo_din_d3[1]_net_1\, 
        \rx_crc_data_store[2]_net_1\, 
        \un1_rx_fifo_din_d3[2]_net_1\, 
        \rx_crc_data_store[3]_net_1\, 
        \un1_rx_fifo_din_d3[3]_net_1\, 
        \rx_crc_data_store[4]_net_1\, 
        \un1_rx_fifo_din_d3[4]_net_1\, 
        \rx_crc_data_store[5]_net_1\, 
        \un1_rx_fifo_din_d3[5]_net_1\, 
        \rx_crc_data_store[6]_net_1\, 
        \un1_rx_fifo_din_d3[6]_net_1\, 
        \rx_crc_data_store[7]_net_1\, 
        \un1_rx_fifo_din_d3[7]_net_1\, 
        \rx_crc_data_store[8]_net_1\, \RX_FIFO_DIN_pipe[0]\, 
        \rx_packet_length[0]_net_1\, N_336_i, 
        \rx_packet_length[1]_net_1\, N_117_i, 
        \rx_packet_length[2]_net_1\, N_119_i, 
        \rx_packet_length[3]_net_1\, 
        \rx_packet_length_13[3]_net_1\, 
        \rx_packet_length[4]_net_1\, 
        \rx_packet_length_13[4]_net_1\, rx_crc_HighByte_en_net_1, 
        ReadFIFO_WR_STATE_1_sqmuxa_1, 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, \RX_FIFO_DIN_pipe[8]\, 
        \ReadFIFO_WR_STATE[3]_net_1\, \rx_end_rst\, N_244_i, 
        N_338_i, N_589, \irx_packet_end\, N_577_i, \RX_EarlyTerm\, 
        \ReadFIFO_WR_STATE[4]_net_1\, \RX_InProcess\, N_311, 
        iRX_FIFO_wr_en_net_1, un5_packet_avail, N_265, 
        \SM_advance_i\, un2_packet_avail, 
        \rx_fifo_din_d2[4]_net_1\, \rx_fifo_din_d1[4]_net_1\, 
        N_236_i, \rx_fifo_din_d2[3]_net_1\, 
        \rx_fifo_din_d1[3]_net_1\, \rx_fifo_din_d2[2]_net_1\, 
        \rx_fifo_din_d1[2]_net_1\, \rx_fifo_din_d2[1]_net_1\, 
        \rx_fifo_din_d1[1]_net_1\, \rx_fifo_din_d2[0]_net_1\, 
        \rx_fifo_din_d1[0]_net_1\, \rx_crc_gen\, 
        un1_ReadFIFO_WR_STATE_15, \rx_fifo_din_d2[7]_net_1\, 
        \rx_fifo_din_d1[7]_net_1\, \rx_fifo_din_d2[6]_net_1\, 
        \rx_fifo_din_d1[6]_net_1\, \rx_fifo_din_d2[5]_net_1\, 
        \rx_fifo_din_d1[5]_net_1\, \ReadFIFO_WR_STATE[8]_net_1\, 
        \ReadFIFO_WR_STATE_ns[1]\, \ReadFIFO_WR_STATE[7]_net_1\, 
        \ReadFIFO_WR_STATE_ns[2]\, \ReadFIFO_WR_STATE[6]_net_1\, 
        \ReadFIFO_WR_STATE_ns[3]\, \ReadFIFO_WR_STATE[5]_net_1\, 
        \ReadFIFO_WR_STATE_ns[4]\, N_225_i, 
        \ReadFIFO_WR_STATE_ns[6]\, \ReadFIFO_WR_STATE[2]_net_1\, 
        \ReadFIFO_WR_STATE_ns[7]\, \ReadFIFO_WR_STATE[1]_net_1\, 
        \ReadFIFO_WR_STATE_ns[8]\, \ReadFIFO_WR_STATE[0]_net_1\, 
        \ReadFIFO_WR_STATE_ns[9]\, \ReadFIFO_WR_STATE[9]_net_1\, 
        N_219_i, RX_InProcess_d1_net_1, \hold_collision\, 
        \N_447_i_i\, un1_tx_collision_detect, 
        \rx_byte_cntr[0]_net_1\, \rx_byte_cntr_s[0]\, N_334_i, 
        \rx_byte_cntr[1]_net_1\, \rx_byte_cntr_s[1]\, 
        \rx_byte_cntr[2]_net_1\, \rx_byte_cntr_s[2]\, 
        \rx_byte_cntr[3]_net_1\, \rx_byte_cntr_s[3]\, 
        \rx_byte_cntr[4]_net_1\, \rx_byte_cntr_s[4]\, 
        \rx_byte_cntr[5]_net_1\, \rx_byte_cntr_s[5]\, 
        \rx_byte_cntr[6]_net_1\, \rx_byte_cntr_s[6]\, 
        \rx_byte_cntr[7]_net_1\, \rx_byte_cntr_s[7]\, 
        \rx_byte_cntr[8]_net_1\, \rx_byte_cntr_s[8]\, 
        \rx_byte_cntr[9]_net_1\, \rx_byte_cntr_s[9]\, 
        \rx_byte_cntr[10]_net_1\, \rx_byte_cntr_s[10]\, 
        \rx_byte_cntr[11]_net_1\, \rx_byte_cntr_s[11]\, 
        rx_byte_cntr_cry_cy, \ReadFIFO_WR_STATE_RNIHSM21_Y[9]\, 
        N_581, \rx_byte_cntr_cry[0]\, \rx_byte_cntr_cry[1]\, 
        \rx_byte_cntr_cry[2]\, \rx_byte_cntr_cry[3]\, 
        \rx_byte_cntr_cry[4]\, \rx_byte_cntr_cry[5]\, 
        \rx_byte_cntr_cry[6]\, \rx_byte_cntr_cry[7]\, 
        \rx_byte_cntr_cry[8]\, \rx_byte_cntr_cry[9]\, 
        \rx_byte_cntr_cry[10]\, \un65_sm_advance_i_cry_0\, 
        \un65_sm_advance_i_cry_1\, un65_sm_advance_i_cry_1_S, 
        \un65_sm_advance_i_cry_2\, un65_sm_advance_i_cry_2_S, 
        \un65_sm_advance_i_cry_3\, un65_sm_advance_i_cry_3_S, 
        \un65_sm_advance_i_cry_4\, un65_sm_advance_i_cry_4_S, 
        \un65_sm_advance_i_cry_5\, un65_sm_advance_i_cry_5_S, 
        \un65_sm_advance_i_cry_6\, un65_sm_advance_i_cry_6_S, 
        \un65_sm_advance_i_cry_7\, un65_sm_advance_i_cry_7_S, 
        \un65_sm_advance_i_cry_8\, un65_sm_advance_i_cry_8_S, 
        \un65_sm_advance_i_cry_9\, un65_sm_advance_i_cry_9_S, 
        \un56_sm_advance_i_cry_0\, \un56_sm_advance_i_cry_1\, 
        un56_sm_advance_i_cry_1_S, \un56_sm_advance_i_cry_2\, 
        un56_sm_advance_i_cry_2_S, \un56_sm_advance_i_cry_3\, 
        un56_sm_advance_i_cry_3_S, \un56_sm_advance_i_cry_4\, 
        un56_sm_advance_i_cry_4_S, \un56_sm_advance_i_cry_5\, 
        un56_sm_advance_i_cry_5_S, \un56_sm_advance_i_cry_6\, 
        un56_sm_advance_i_cry_6_S, \un56_sm_advance_i_cry_7\, 
        un56_sm_advance_i_cry_7_S, \un56_sm_advance_i_cry_8\, 
        un56_sm_advance_i_cry_8_S, \un56_sm_advance_i_cry_9\, 
        un56_sm_advance_i_cry_9_S, un67_sm_advance_i_cry_0, 
        un67_sm_advance_i_cry_1, un67_sm_advance_i_cry_2, 
        un67_sm_advance_i_cry_3, un67_sm_advance_i_cry_4, 
        un67_sm_advance_i_cry_5, un67_sm_advance_i_cry_6, 
        un67_sm_advance_i_cry_7, un67_sm_advance_i_cry_8, 
        un67_sm_advance_i_cry_9, un67_sm_advance_i_cry_10, 
        un67_sm_advance_i, \un58_sm_advance_i_0_data_tmp[0]\, 
        \un58_sm_advance_i_0_data_tmp[1]\, 
        \un58_sm_advance_i_0_data_tmp[2]\, 
        \un58_sm_advance_i_0_data_tmp[3]\, 
        \un58_sm_advance_i_0_data_tmp[4]\, 
        \un58_sm_advance_i_0_data_tmp[5]\, 
        \un1_sampler_clk1x_en_0_data_tmp[0]\, 
        \rx_crc_data_calc[0]\, \rx_crc_data_calc[1]\, 
        \un1_sampler_clk1x_en_0_data_tmp[1]\, 
        \rx_crc_data_calc[2]\, \rx_crc_data_calc[3]\, 
        \un1_sampler_clk1x_en_0_data_tmp[2]\, 
        \rx_crc_data_calc[4]\, \rx_crc_data_calc[5]\, 
        \un1_sampler_clk1x_en_0_data_tmp[3]\, 
        \rx_crc_data_calc[6]\, \rx_crc_data_calc[7]\, 
        \un1_sampler_clk1x_en_0_data_tmp[4]\, 
        \rx_crc_data_calc[8]\, \rx_crc_data_calc[9]\, 
        \un1_sampler_clk1x_en_0_data_tmp[5]\, 
        \rx_crc_data_calc[10]\, \rx_crc_data_calc[11]\, 
        \un1_sampler_clk1x_en_0_data_tmp[6]\, 
        \rx_crc_data_calc[12]\, \rx_crc_data_calc[13]\, 
        \un1_sampler_clk1x_en_0_data_tmp[7]\, 
        \rx_crc_data_calc[14]\, \rx_crc_data_calc[15]\, N_97, 
        \ReadFIFO_WR_STATE_ns_i_0_a2_3_0[5]_net_1\, 
        \ReadFIFO_WR_STATE_ns_i_0_a2_d[5]_net_1\, N_225_i_1, 
        \ReadFIFO_WR_STATE_ns_i_0_a2_0_0[5]_net_1\, 
        un40_sm_advance_i_1, un40_sm_advance_i_2, 
        \ReadFIFO_WR_STATE_ns_0_a2_0_1_1[3]_net_1\, 
        un1_ReadFIFO_WR_STATE_14_0_0_a2_0, un38_sm_advance_i_3, 
        un35_sm_advance_i_3, un32_sm_advance_i_3, 
        un29_sm_advance_i_7, N_582, N_269, N_282, 
        consumer_type_12_sn_N_2, rx_byte_cntrlde_i_a2_0_0, 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0_a2_0\, 
        un29_sm_advance_i_NE_4, un29_sm_advance_i_NE_3, 
        un29_sm_advance_i_NE_2, un29_sm_advance_i_NE_1, 
        un32_sm_advance_i_NE_4, un32_sm_advance_i_NE_3, 
        un32_sm_advance_i_NE_1, un32_sm_advance_i_NE_0, 
        un35_sm_advance_i_NE_4, un35_sm_advance_i_NE_3, 
        un35_sm_advance_i_NE_1, un35_sm_advance_i_NE_0, 
        un38_sm_advance_i_NE_4, un38_sm_advance_i_NE_3, 
        un38_sm_advance_i_NE_1, un38_sm_advance_i_NE_0, N_275, 
        N_670, N_294, N_273, 
        \ReadFIFO_WR_STATE_ns_0_a2_0_0[6]_net_1\, 
        un29_sm_advance_i_NE_5, un32_sm_advance_i_NE_6, 
        un35_sm_advance_i_NE_6, un38_sm_advance_i_NE_6, N_405, 
        N_417, N_396, \ReadFIFO_WR_STATE_ns_0_0[4]_net_1\, 
        un32_sm_advance_i_NE_7, un35_sm_advance_i_NE_7, 
        un38_sm_advance_i_NE_7, un30_sm_advance_i : std_logic;

    for all : CRC16_Generator_1
	Use entity work.CRC16_Generator_1(DEF_ARCH);
begin 

    RX_FIFO_DIN_pipe(8) <= \RX_FIFO_DIN_pipe[8]\;
    RX_FIFO_DIN_pipe(7) <= \RX_FIFO_DIN_pipe[7]\;
    RX_FIFO_DIN_pipe(6) <= \RX_FIFO_DIN_pipe[6]\;
    RX_FIFO_DIN_pipe(5) <= \RX_FIFO_DIN_pipe[5]\;
    RX_FIFO_DIN_pipe(4) <= \RX_FIFO_DIN_pipe[4]\;
    RX_FIFO_DIN_pipe(3) <= \RX_FIFO_DIN_pipe[3]\;
    RX_FIFO_DIN_pipe(2) <= \RX_FIFO_DIN_pipe[2]\;
    RX_FIFO_DIN_pipe(1) <= \RX_FIFO_DIN_pipe[1]\;
    RX_FIFO_DIN_pipe(0) <= \RX_FIFO_DIN_pipe[0]\;
    N_447_i_i <= \N_447_i_i\;
    RX_InProcess_d1 <= RX_InProcess_d1_net_1;
    iRX_FIFO_wr_en <= iRX_FIFO_wr_en_net_1;
    RX_EarlyTerm <= \RX_EarlyTerm\;
    rx_crc_HighByte_en <= rx_crc_HighByte_en_net_1;
    rx_packet_complt <= rx_packet_complt_net_1;
    rx_CRC_error <= rx_CRC_error_net_1;

    un56_sm_advance_i_cry_8 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[9]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un56_sm_advance_i_cry_7\, S => un56_sm_advance_i_cry_8_S, 
        Y => OPEN, FCO => \un56_sm_advance_i_cry_8\);
    
    \rx_packet_length[5]\ : SLE
      port map(D => \rx_packet_length_13[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \un1_ReadFIFO_WR_STATE_14_0_0\, 
        ALn => N_480_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[5]_net_1\);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE_7\ : CFG3
      generic map(INIT => x"FE")

      port map(A => un32_sm_advance_i_NE_4, B => 
        un32_sm_advance_i_NE_1, C => un32_sm_advance_i_NE_0, Y
         => un32_sm_advance_i_NE_7);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_4\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type3_reg(9), B => 
        consumer_type3_reg(2), C => \consumer_type[9]_net_1\, D
         => \consumer_type[2]_net_1\, Y => un35_sm_advance_i_NE_4);
    
    \ReadFIFO_WRITE_PROC.un5_packet_avail_0_a2\ : CFG3
      generic map(INIT => x"80")

      port map(A => \bit_cntr[2]_net_1\, B => \bit_cntr[1]_net_1\, 
        C => \bit_cntr[0]_net_1\, Y => un5_packet_avail);
    
    \rx_packet_length_RNO[1]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => N_282, B => N_273, C => 
        \rx_packet_length[1]_net_1\, D => RX_FIFO_DIN(1), Y => 
        N_117_i);
    
    N_447_i : CFG2
      generic map(INIT => x"1")

      port map(A => idle_line, B => N_480, Y => \N_447_i_i\);
    
    consumer_type_0_sqmuxa_0_a3_i : CFG3
      generic map(INIT => x"80")

      port map(A => packet_avail, B => 
        \ReadFIFO_WR_STATE[9]_net_1\, C => N_236_i, Y => N_97);
    
    rx_crc_LowByte_en : SLE
      port map(D => \ReadFIFO_WR_STATE[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[8]\);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE_7\ : CFG3
      generic map(INIT => x"FE")

      port map(A => un38_sm_advance_i_NE_4, B => 
        un38_sm_advance_i_NE_1, C => un38_sm_advance_i_NE_0, Y
         => un38_sm_advance_i_NE_7);
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_27\ : ARI1
      generic map(INIT => x"68241")

      port map(A => un56_sm_advance_i_cry_7_S, B => 
        \rx_byte_cntr[8]_net_1\, C => \rx_byte_cntr[9]_net_1\, D
         => un56_sm_advance_i_cry_8_S, FCI => 
        \un58_sm_advance_i_0_data_tmp[3]\, S => OPEN, Y => OPEN, 
        FCO => \un58_sm_advance_i_0_data_tmp[4]\);
    
    un56_sm_advance_i_cry_6 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[7]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un56_sm_advance_i_cry_5\, S => un56_sm_advance_i_cry_6_S, 
        Y => OPEN, FCO => \un56_sm_advance_i_cry_6\);
    
    \SM_advancebit_cntr_RNO[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => N_265, B => \SM_advancebit_cntr[0]_net_1\, Y
         => N_321_i_i);
    
    \rx_packet_length[10]\ : SLE
      port map(D => N_125_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_ReadFIFO_WR_STATE_14_0_0\, ALn => N_480_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_packet_length[10]_net_1\);
    
    un1_ReadFIFO_WR_STATE_15_0_a2 : CFG4
      generic map(INIT => x"0400")

      port map(A => \hold_collision\, B => 
        \ReadFIFO_WR_STATE[5]_net_1\, C => un67_sm_advance_i, D
         => \un58_sm_advance_i_0_data_tmp[5]\, Y => N_417);
    
    un1_iRX_EarlyTerm_1_sqmuxa_1_0_0 : CFG4
      generic map(INIT => x"F1F0")

      port map(A => \ReadFIFO_WR_STATE[8]_net_1\, B => N_311, C
         => N_236_i, D => \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0_a2_0\, 
        Y => \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\);
    
    \rx_byte_cntr[11]\ : SLE
      port map(D => \rx_byte_cntr_s[11]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_334_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_byte_cntr[11]_net_1\);
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_33\ : ARI1
      generic map(INIT => x"68241")

      port map(A => un56_sm_advance_i_cry_3_S, B => 
        \rx_byte_cntr[4]_net_1\, C => \rx_byte_cntr[5]_net_1\, D
         => un56_sm_advance_i_cry_4_S, FCI => 
        \un58_sm_advance_i_0_data_tmp[1]\, S => OPEN, Y => OPEN, 
        FCO => \un58_sm_advance_i_0_data_tmp[2]\);
    
    \ReadFIFO_WR_STATE[4]\ : SLE
      port map(D => N_225_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_WR_STATE[4]_net_1\);
    
    \rx_byte_cntr_RNIT3CF2[0]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \rx_byte_cntr[0]_net_1\, C
         => \ReadFIFO_WR_STATE_RNIHSM21_Y[9]\, D => GND_net_1, 
        FCI => rx_byte_cntr_cry_cy, S => \rx_byte_cntr_s[0]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[0]\);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE_2\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type1_reg(4), B => 
        consumer_type1_reg(3), C => \consumer_type[4]_net_1\, D
         => \consumer_type[3]_net_1\, Y => un29_sm_advance_i_NE_2);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_6\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[6]_net_1\, B => 
        un65_sm_advance_i_cry_5_S, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_5, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_6);
    
    rx_end_rst : SLE
      port map(D => N_244_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => N_480_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_end_rst\);
    
    \ReadFIFO_WR_STATE_ns_i_0_a2_d[5]\ : CFG4
      generic map(INIT => x"0111")

      port map(A => \ReadFIFO_WR_STATE[4]_net_1\, B => 
        \hold_collision\, C => un40_sm_advance_i_2, D => 
        un40_sm_advance_i_1, Y => 
        \ReadFIFO_WR_STATE_ns_i_0_a2_d[5]_net_1\);
    
    un1_ReadFIFO_WR_STATE_14_0_0_o2_RNIDF0U : CFG4
      generic map(INIT => x"5100")

      port map(A => N_311, B => \ReadFIFO_WR_STATE[2]_net_1\, C
         => N_236_i, D => N_269, Y => N_333_i);
    
    \ReadFIFO_WR_STATE_ns_0[6]\ : CFG4
      generic map(INIT => x"22F2")

      port map(A => \ReadFIFO_WR_STATE[3]_net_1\, B => N_236_i, C
         => \ReadFIFO_WR_STATE_ns_0_a2_0_0[6]_net_1\, D => 
        \un58_sm_advance_i_0_data_tmp[5]\, Y => 
        \ReadFIFO_WR_STATE_ns[6]\);
    
    \rx_fifo_din_d3[2]\ : SLE
      port map(D => \rx_fifo_din_d2[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_236_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[2]\);
    
    \SM_advancebit_cntr[0]\ : SLE
      port map(D => N_321_i_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un8_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SM_advancebit_cntr[0]_net_1\);
    
    \iRX_FIFO_wr_en\ : SLE
      port map(D => un5_packet_avail, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_265, ALn => un15_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        iRX_FIFO_wr_en_net_1);
    
    \rx_packet_length[8]\ : SLE
      port map(D => N_337_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_ReadFIFO_WR_STATE_14_0_0\, ALn => N_480_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_packet_length[8]_net_1\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_1\ : ARI1
      generic map(INIT => x"555AA")

      port map(A => \rx_byte_cntr[1]_net_1\, B => 
        \rx_packet_length[1]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => un67_sm_advance_i_cry_0, S => OPEN, Y
         => OPEN, FCO => un67_sm_advance_i_cry_1);
    
    \consumer_type[4]\ : SLE
      port map(D => \consumer_type_12[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_333_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type[4]_net_1\);
    
    \rx_fifo_din_d1[0]\ : SLE
      port map(D => RX_FIFO_DIN(0), CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_236_i, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_fifo_din_d1[0]_net_1\);
    
    \ReadFIFO_WR_STATE_ns_0_a2_0_1_1[3]\ : CFG4
      generic map(INIT => x"440F")

      port map(A => \hold_collision\, B => 
        \ReadFIFO_WR_STATE[7]_net_1\, C => 
        \ReadFIFO_WR_STATE[6]_net_1\, D => N_236_i, Y => 
        \ReadFIFO_WR_STATE_ns_0_a2_0_1_1[3]_net_1\);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE_0\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type4_reg(8), B => 
        consumer_type4_reg(7), C => \consumer_type[8]_net_1\, D
         => \consumer_type[7]_net_1\, Y => un38_sm_advance_i_NE_0);
    
    \rx_crc_data_store[1]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_330_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_store[1]_net_1\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_11\ : ARI1
      generic map(INIT => x"555AA")

      port map(A => \rx_byte_cntr[11]_net_1\, B => 
        \un65_sm_advance_i_cry_9\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_10, S => OPEN, Y => OPEN, 
        FCO => un67_sm_advance_i);
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_9\ : ARI1
      generic map(INIT => x"62184")

      port map(A => \un56_sm_advance_i_cry_9\, B => 
        \rx_byte_cntr[10]_net_1\, C => \rx_byte_cntr[11]_net_1\, 
        D => un56_sm_advance_i_cry_9_S, FCI => 
        \un58_sm_advance_i_0_data_tmp[4]\, S => OPEN, Y => OPEN, 
        FCO => \un58_sm_advance_i_0_data_tmp[5]\);
    
    \un1_rx_fifo_din_d3[4]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[4]\, B => 
        rx_crc_HighByte_en_net_1, Y => 
        \un1_rx_fifo_din_d3[4]_net_1\);
    
    un1_ReadFIFO_WR_STATE_7_i_a3_i_o2 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \ReadFIFO_WR_STATE[7]_net_1\, B => 
        \ReadFIFO_WR_STATE[6]_net_1\, C => 
        \ReadFIFO_WR_STATE[5]_net_1\, D => 
        \ReadFIFO_WR_STATE[3]_net_1\, Y => N_311);
    
    \rx_fifo_din_d3[4]\ : SLE
      port map(D => \rx_fifo_din_d2[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_236_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[4]\);
    
    \consumer_type[7]\ : SLE
      port map(D => \consumer_type_12[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_333_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type[7]_net_1\);
    
    \ReadFIFO_WR_STATE_RNO[9]\ : CFG4
      generic map(INIT => x"0CEE")

      port map(A => idle_line, B => \ReadFIFO_WR_STATE[9]_net_1\, 
        C => N_97, D => N_582, Y => N_219_i);
    
    \rx_byte_cntr_RNI14NKD[8]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \rx_byte_cntr[8]_net_1\, C
         => \ReadFIFO_WR_STATE_RNIHSM21_Y[9]\, D => GND_net_1, 
        FCI => \rx_byte_cntr_cry[7]\, S => \rx_byte_cntr_s[8]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[8]\);
    
    \ReadFIFO_WR_SM.consumer_type_12[9]\ : CFG4
      generic map(INIT => x"CCA0")

      port map(A => RX_FIFO_DIN(7), B => \consumer_type[9]_net_1\, 
        C => N_97, D => \ReadFIFO_WR_STATE[8]_net_1\, Y => 
        \consumer_type_12[9]\);
    
    un65_sm_advance_i_cry_2 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[3]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un65_sm_advance_i_cry_1\, S => un65_sm_advance_i_cry_2_S, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_2\);
    
    \rx_fifo_din_d1[5]\ : SLE
      port map(D => RX_FIFO_DIN(5), CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_236_i, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_fifo_din_d1[5]_net_1\);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_45\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[9]_net_1\, B => 
        \rx_crc_data_calc[8]\, C => \rx_crc_data_calc[9]\, D => 
        \rx_crc_data_store[8]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[3]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[4]\);
    
    \rx_crc_data_store[12]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_344_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_store[12]_net_1\);
    
    \rx_crc_HighByte_en\ : SLE
      port map(D => ReadFIFO_WR_STATE_1_sqmuxa_1, CLK => 
        CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rx_crc_HighByte_en_net_1);
    
    un56_sm_advance_i_cry_1 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[2]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un56_sm_advance_i_cry_0\, S => un56_sm_advance_i_cry_1_S, 
        Y => OPEN, FCO => \un56_sm_advance_i_cry_1\);
    
    \HOLD_COL_PROC.un1_tx_collision_detect\ : CFG2
      generic map(INIT => x"8")

      port map(A => TX_collision_detect, B => tx_col_detect_en, Y
         => un1_tx_collision_detect);
    
    \rx_CRC_error\ : SLE
      port map(D => N_589, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rx_CRC_error_net_1);
    
    \rx_crc_data_store[8]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_344_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_store[8]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \rx_byte_cntr_RNIOLM85[2]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \rx_byte_cntr[2]_net_1\, C
         => \ReadFIFO_WR_STATE_RNIHSM21_Y[9]\, D => GND_net_1, 
        FCI => \rx_byte_cntr_cry[1]\, S => \rx_byte_cntr_s[2]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[2]\);
    
    \rx_fifo_din_d1[2]\ : SLE
      port map(D => RX_FIFO_DIN(2), CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_236_i, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_fifo_din_d1[2]_net_1\);
    
    \consumer_type[6]\ : SLE
      port map(D => \consumer_type_12[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_333_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type[6]_net_1\);
    
    \rx_crc_data_store[5]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_330_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_store[5]_net_1\);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_9\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[3]_net_1\, B => 
        \rx_crc_data_calc[2]\, C => \rx_crc_data_calc[3]\, D => 
        \rx_crc_data_store[2]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[0]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[1]\);
    
    \rx_byte_cntr_RNIJDCCG[10]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \rx_byte_cntr[10]_net_1\, C
         => \ReadFIFO_WR_STATE_RNIHSM21_Y[9]\, D => GND_net_1, 
        FCI => \rx_byte_cntr_cry[9]\, S => \rx_byte_cntr_s[10]\, 
        Y => OPEN, FCO => \rx_byte_cntr_cry[10]\);
    
    \rx_packet_length[6]\ : SLE
      port map(D => \rx_packet_length_13[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \un1_ReadFIFO_WR_STATE_14_0_0\, 
        ALn => N_480_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[6]_net_1\);
    
    \ReadFIFO_WR_STATE[2]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \ReadFIFO_WR_STATE[2]_net_1\);
    
    \rx_byte_cntr[1]\ : SLE
      port map(D => \rx_byte_cntr_s[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_334_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_byte_cntr[1]_net_1\);
    
    \ReadFIFO_WR_STATE_RNIHSM21[9]\ : ARI1
      generic map(INIT => x"4B300")

      port map(A => N_581, B => N_236_i, C => 
        \ReadFIFO_WR_STATE[9]_net_1\, D => packet_avail, FCI => 
        VCC_net_1, S => OPEN, Y => 
        \ReadFIFO_WR_STATE_RNIHSM21_Y[9]\, FCO => 
        rx_byte_cntr_cry_cy);
    
    un56_sm_advance_i_cry_4 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[5]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un56_sm_advance_i_cry_3\, S => un56_sm_advance_i_cry_4_S, 
        Y => OPEN, FCO => \un56_sm_advance_i_cry_4\);
    
    \rx_packet_length_13_i_o2[8]\ : CFG2
      generic map(INIT => x"D")

      port map(A => N_236_i, B => \ReadFIFO_WR_STATE[6]_net_1\, Y
         => N_275);
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_1\ : ARI1
      generic map(INIT => x"62184")

      port map(A => \rx_packet_length[1]_net_1\, B => 
        \rx_byte_cntr[0]_net_1\, C => \rx_byte_cntr[1]_net_1\, D
         => \rx_packet_length[0]_net_1\, FCI => GND_net_1, S => 
        OPEN, Y => OPEN, FCO => \un58_sm_advance_i_0_data_tmp[0]\);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE_1\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type4_reg(6), B => 
        consumer_type4_reg(5), C => \consumer_type[6]_net_1\, D
         => \consumer_type[5]_net_1\, Y => un38_sm_advance_i_NE_1);
    
    un65_sm_advance_i_cry_6 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[7]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un65_sm_advance_i_cry_5\, S => un65_sm_advance_i_cry_6_S, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_6\);
    
    \ReadFIFO_WR_STATE_ns_0_a2_0[1]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => packet_avail, B => \hold_collision\, C => 
        N_236_i, D => \ReadFIFO_WR_STATE[9]_net_1\, Y => N_396);
    
    \rx_packet_complt\ : SLE
      port map(D => N_338_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rx_packet_complt_net_1);
    
    iRX_EarlyTerm : SLE
      port map(D => \ReadFIFO_WR_STATE[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_EarlyTerm\);
    
    \ReadFIFO_WR_SM.consumer_type_12[4]\ : CFG4
      generic map(INIT => x"F088")

      port map(A => RX_FIFO_DIN(2), B => N_97, C => 
        \consumer_type[4]_net_1\, D => 
        \ReadFIFO_WR_STATE[8]_net_1\, Y => \consumer_type_12[4]\);
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_21\ : ARI1
      generic map(INIT => x"68241")

      port map(A => un56_sm_advance_i_cry_5_S, B => 
        \rx_byte_cntr[6]_net_1\, C => \rx_byte_cntr[7]_net_1\, D
         => un56_sm_advance_i_cry_6_S, FCI => 
        \un58_sm_advance_i_0_data_tmp[2]\, S => OPEN, Y => OPEN, 
        FCO => \un58_sm_advance_i_0_data_tmp[3]\);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE_4\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type4_reg(9), B => 
        consumer_type4_reg(2), C => \consumer_type[9]_net_1\, D
         => \consumer_type[2]_net_1\, Y => un38_sm_advance_i_NE_4);
    
    un65_sm_advance_i_cry_3 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[4]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un65_sm_advance_i_cry_2\, S => un65_sm_advance_i_cry_3_S, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_3\);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_21\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[15]_net_1\, B => 
        \rx_crc_data_calc[14]\, C => \rx_crc_data_calc[15]\, D
         => \rx_crc_data_store[14]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[6]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[7]\);
    
    \ReadFIFO_WR_STATE_ns_i_0_a2_0_0[5]\ : CFG3
      generic map(INIT => x"07")

      port map(A => packet_avail, B => 
        \ReadFIFO_WR_STATE[9]_net_1\, C => 
        \ReadFIFO_WR_STATE[4]_net_1\, Y => 
        \ReadFIFO_WR_STATE_ns_i_0_a2_0_0[5]_net_1\);
    
    \bit_cntr[2]\ : SLE
      port map(D => N_350_i_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un15_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \bit_cntr[2]_net_1\);
    
    rx_packet_complt_RNO : CFG3
      generic map(INIT => x"20")

      port map(A => idle_line, B => tx_col_detect_en, C => 
        \ReadFIFO_WR_STATE[0]_net_1\, Y => N_338_i);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => un29_sm_advance_i_NE_2, B => 
        un29_sm_advance_i_NE_5, C => un29_sm_advance_i_NE_4, D
         => un29_sm_advance_i_NE_3, Y => un30_sm_advance_i);
    
    \rx_packet_length_13[3]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => N_282, B => N_273, C => 
        \rx_packet_length[3]_net_1\, D => RX_FIFO_DIN(3), Y => 
        \rx_packet_length_13[3]_net_1\);
    
    \bit_cntr[0]\ : SLE
      port map(D => N_322_i_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un15_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \bit_cntr[0]_net_1\);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE_4\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type1_reg(9), B => 
        consumer_type1_reg(2), C => \consumer_type[9]_net_1\, D
         => \consumer_type[2]_net_1\, Y => un29_sm_advance_i_NE_4);
    
    un56_sm_advance_i_cry_9 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[10]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un56_sm_advance_i_cry_8\, S => un56_sm_advance_i_cry_9_S, 
        Y => OPEN, FCO => \un56_sm_advance_i_cry_9\);
    
    un56_sm_advance_i_cry_3 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[4]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un56_sm_advance_i_cry_2\, S => un56_sm_advance_i_cry_3_S, 
        Y => OPEN, FCO => \un56_sm_advance_i_cry_3\);
    
    \rx_packet_length_13[5]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => N_282, B => N_273, C => 
        \rx_packet_length[5]_net_1\, D => RX_FIFO_DIN(5), Y => 
        \rx_packet_length_13[5]_net_1\);
    
    \rx_packet_length_13[6]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => N_282, B => N_273, C => 
        \rx_packet_length[6]_net_1\, D => RX_FIFO_DIN(6), Y => 
        \rx_packet_length_13[6]_net_1\);
    
    un1_ReadFIFO_WR_STATE_14_0_0 : CFG4
      generic map(INIT => x"CCCE")

      port map(A => N_236_i, B => N_405, C => 
        \ReadFIFO_WR_STATE[5]_net_1\, D => 
        \ReadFIFO_WR_STATE[3]_net_1\, Y => 
        \un1_ReadFIFO_WR_STATE_14_0_0\);
    
    un1_ReadFIFO_WR_STATE_15_0_0 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \ReadFIFO_WR_STATE[8]_net_1\, B => 
        \ReadFIFO_WR_STATE[9]_net_1\, C => N_417, D => N_282, Y
         => un1_ReadFIFO_WR_STATE_15);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \ReadFIFO_WR_STATE[7]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \ReadFIFO_WR_STATE[7]_net_1\);
    
    \rx_fifo_din_d2[6]\ : SLE
      port map(D => \rx_fifo_din_d1[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_236_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_fifo_din_d2[6]_net_1\);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE_6\ : CFG4
      generic map(INIT => x"FFF6")

      port map(A => \consumer_type[4]_net_1\, B => 
        consumer_type2_reg(4), C => un32_sm_advance_i_NE_3, D => 
        un32_sm_advance_i_3, Y => un32_sm_advance_i_NE_6);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE_6\ : CFG4
      generic map(INIT => x"FFF6")

      port map(A => \consumer_type[4]_net_1\, B => 
        consumer_type4_reg(4), C => un38_sm_advance_i_NE_3, D => 
        un38_sm_advance_i_3, Y => un38_sm_advance_i_NE_6);
    
    \rx_packet_length[2]\ : SLE
      port map(D => N_119_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_ReadFIFO_WR_STATE_14_0_0\, ALn => N_480_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_packet_length[2]_net_1\);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_3\ : CFG2
      generic map(INIT => x"6")

      port map(A => \consumer_type[3]_net_1\, B => 
        consumer_type3_reg(3), Y => un35_sm_advance_i_3);
    
    \rx_fifo_din_d2[0]\ : SLE
      port map(D => \rx_fifo_din_d1[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_236_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_fifo_din_d2[0]_net_1\);
    
    \ReadFIFO_WR_STATE_RNO[4]\ : CFG4
      generic map(INIT => x"1011")

      port map(A => \ReadFIFO_WR_STATE_ns_i_0_a2_3_0[5]_net_1\, B
         => \ReadFIFO_WR_STATE_ns_i_0_a2_d[5]_net_1\, C => N_311, 
        D => N_225_i_1, Y => N_225_i);
    
    \ReadFIFO_WR_STATE_RNI3DOS1[9]\ : CFG4
      generic map(INIT => x"23AF")

      port map(A => \ReadFIFO_WR_STATE[9]_net_1\, B => 
        rx_byte_cntrlde_i_a2_0_0, C => N_294, D => 
        \ReadFIFO_WR_STATE_RNIHSM21_Y[9]\, Y => N_334_i);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_8\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[8]_net_1\, B => 
        un65_sm_advance_i_cry_7_S, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_7, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_8);
    
    \SM_advancebit_cntr[1]\ : SLE
      port map(D => N_325_i_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un8_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SM_advancebit_cntr[1]_net_1\);
    
    \bit_cntr[1]\ : SLE
      port map(D => N_326_i_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un15_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \bit_cntr[1]_net_1\);
    
    \rx_byte_cntr[9]\ : SLE
      port map(D => \rx_byte_cntr_s[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_334_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_byte_cntr[9]_net_1\);
    
    \un1_rx_fifo_din_d3[1]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[1]\, B => 
        rx_crc_HighByte_en_net_1, Y => 
        \un1_rx_fifo_din_d3[1]_net_1\);
    
    \rx_crc_data_store[13]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_344_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_store[13]_net_1\);
    
    \rx_crc_data_store[0]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_330_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_store[0]_net_1\);
    
    \rx_byte_cntr_RNIAC1S3[1]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \rx_byte_cntr[1]_net_1\, C
         => \ReadFIFO_WR_STATE_RNIHSM21_Y[9]\, D => GND_net_1, 
        FCI => \rx_byte_cntr_cry[0]\, S => \rx_byte_cntr_s[1]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[1]\);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_15\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[5]_net_1\, B => 
        \rx_crc_data_calc[4]\, C => \rx_crc_data_calc[5]\, D => 
        \rx_crc_data_store[4]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[1]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[2]\);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_0\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type3_reg(8), B => 
        consumer_type3_reg(7), C => \consumer_type[8]_net_1\, D
         => \consumer_type[7]_net_1\, Y => un35_sm_advance_i_NE_0);
    
    \ReadFIFO_WR_STATE_ns_0[8]\ : CFG3
      generic map(INIT => x"D5")

      port map(A => N_269, B => N_236_i, C => 
        \ReadFIFO_WR_STATE[2]_net_1\, Y => 
        \ReadFIFO_WR_STATE_ns[8]\);
    
    \consumer_type[1]\ : SLE
      port map(D => \consumer_type_12[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_333_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type[1]_net_1\);
    
    \bit_cntr_RNO[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => N_265, B => \bit_cntr[0]_net_1\, Y => 
        N_322_i_i);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_4\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[4]_net_1\, B => 
        un65_sm_advance_i_cry_3_S, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_3, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_4);
    
    \rx_fifo_din_d1[4]\ : SLE
      port map(D => RX_FIFO_DIN(4), CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_236_i, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_fifo_din_d1[4]_net_1\);
    
    SM_advance_i_RNIR6AL : CFG3
      generic map(INIT => x"37")

      port map(A => \ReadFIFO_WR_STATE[1]_net_1\, B => 
        sampler_clk1x_en, C => \SM_advance_i\, Y => N_294);
    
    \rx_fifo_din_d2[1]\ : SLE
      port map(D => \rx_fifo_din_d1[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_236_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_fifo_din_d2[1]_net_1\);
    
    \rx_packet_length_RNO[10]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => N_282, B => N_275, C => 
        \rx_packet_length[10]_net_1\, D => RX_FIFO_DIN(2), Y => 
        N_125_i);
    
    \un1_rx_fifo_din_d3[7]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[7]\, B => 
        rx_crc_HighByte_en_net_1, Y => 
        \un1_rx_fifo_din_d3[7]_net_1\);
    
    \rx_packet_length_RNO[8]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => N_282, B => N_275, C => 
        \rx_packet_length[8]_net_1\, D => RX_FIFO_DIN(0), Y => 
        N_337_i);
    
    \ReadFIFO_WR_STATE[0]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \ReadFIFO_WR_STATE[0]_net_1\);
    
    \ReadFIFO_WR_STATE[6]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \ReadFIFO_WR_STATE[6]_net_1\);
    
    \rx_fifo_din_d2[5]\ : SLE
      port map(D => \rx_fifo_din_d1[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_236_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_fifo_din_d2[5]_net_1\);
    
    \rx_fifo_din_d1[3]\ : SLE
      port map(D => RX_FIFO_DIN(3), CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_236_i, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_fifo_din_d1[3]_net_1\);
    
    \un1_rx_fifo_din_d3[0]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[0]\, B => 
        rx_crc_HighByte_en_net_1, Y => 
        \un1_rx_fifo_din_d3[0]_net_1\);
    
    \ReadFIFO_WR_STATE_ns_0_a2_0_1[3]\ : CFG4
      generic map(INIT => x"4C33")

      port map(A => un40_sm_advance_i_1, B => N_236_i, C => 
        un40_sm_advance_i_2, D => 
        \ReadFIFO_WR_STATE_ns_0_a2_0_1_1[3]_net_1\, Y => 
        \ReadFIFO_WR_STATE_ns[3]\);
    
    \ReadFIFO_WR_SM.un40_sm_advance_i_1\ : CFG4
      generic map(INIT => x"EEE0")

      port map(A => un38_sm_advance_i_NE_7, B => 
        un38_sm_advance_i_NE_6, C => un35_sm_advance_i_NE_7, D
         => un35_sm_advance_i_NE_6, Y => un40_sm_advance_i_1);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_9\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[9]_net_1\, B => 
        un65_sm_advance_i_cry_8_S, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_8, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_9);
    
    consumer_type_0_sqmuxa_0_a3_i_RNIST29 : CFG2
      generic map(INIT => x"1")

      port map(A => N_97, B => \ReadFIFO_WR_STATE[8]_net_1\, Y
         => consumer_type_12_sn_N_2);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_7\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[7]_net_1\, B => 
        un65_sm_advance_i_cry_6_S, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_6, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_7);
    
    \ReadFIFO_WR_SM.consumer_type_12[6]\ : CFG4
      generic map(INIT => x"F088")

      port map(A => RX_FIFO_DIN(4), B => N_97, C => 
        \consumer_type[6]_net_1\, D => 
        \ReadFIFO_WR_STATE[8]_net_1\, Y => \consumer_type_12[6]\);
    
    \rx_byte_cntr_RNI8OME9[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \rx_byte_cntr[5]_net_1\, C
         => \ReadFIFO_WR_STATE_RNIHSM21_Y[9]\, D => GND_net_1, 
        FCI => \rx_byte_cntr_cry[4]\, S => \rx_byte_cntr_s[5]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[5]\);
    
    \rx_byte_cntr[8]\ : SLE
      port map(D => \rx_byte_cntr_s[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_334_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_byte_cntr[8]_net_1\);
    
    \rx_byte_cntr[2]\ : SLE
      port map(D => \rx_byte_cntr_s[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_334_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_byte_cntr[2]_net_1\);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE_1\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type2_reg(6), B => 
        consumer_type2_reg(5), C => \consumer_type[6]_net_1\, D
         => \consumer_type[5]_net_1\, Y => un32_sm_advance_i_NE_1);
    
    \ReadFIFO_WR_STATE_ns_0_o2[4]\ : CFG2
      generic map(INIT => x"7")

      port map(A => N_236_i, B => \ReadFIFO_WR_STATE[6]_net_1\, Y
         => N_273);
    
    \rx_packet_length_RNO[9]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => N_282, B => N_275, C => 
        \rx_packet_length[9]_net_1\, D => RX_FIFO_DIN(1), Y => 
        N_123_i);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_7\ : CFG3
      generic map(INIT => x"FE")

      port map(A => un35_sm_advance_i_NE_4, B => 
        un35_sm_advance_i_NE_1, C => un35_sm_advance_i_NE_0, Y
         => un35_sm_advance_i_NE_7);
    
    \rx_packet_length[7]\ : SLE
      port map(D => \rx_packet_length_13[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \un1_ReadFIFO_WR_STATE_14_0_0\, 
        ALn => N_480_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[7]_net_1\);
    
    un56_sm_advance_i_cry_0 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[1]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => GND_net_1, S => 
        OPEN, Y => OPEN, FCO => \un56_sm_advance_i_cry_0\);
    
    \SM_ADVANCE_PROC.un2_packet_avail_0_a2\ : CFG3
      generic map(INIT => x"80")

      port map(A => \SM_advancebit_cntr[2]_net_1\, B => 
        \SM_advancebit_cntr[1]_net_1\, C => 
        \SM_advancebit_cntr[0]_net_1\, Y => un2_packet_avail);
    
    \ReadFIFO_WR_SM.consumer_type_12[0]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => RX_FIFO_DIN(6), B => \consumer_type[0]_net_1\, 
        C => consumer_type_12_sn_N_2, D => N_670, Y => 
        \consumer_type_12[0]\);
    
    un1_ReadFIFO_WR_STATE_14_0_0_a2_0_0 : CFG2
      generic map(INIT => x"1")

      port map(A => \ReadFIFO_WR_STATE[8]_net_1\, B => 
        \ReadFIFO_WR_STATE[2]_net_1\, Y => 
        un1_ReadFIFO_WR_STATE_14_0_0_a2_0);
    
    \rx_byte_cntr_RNIQ5CRA[6]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \rx_byte_cntr[6]_net_1\, C
         => \ReadFIFO_WR_STATE_RNIHSM21_Y[9]\, D => GND_net_1, 
        FCI => \rx_byte_cntr_cry[5]\, S => \rx_byte_cntr_s[6]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[6]\);
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_15\ : ARI1
      generic map(INIT => x"68241")

      port map(A => un56_sm_advance_i_cry_1_S, B => 
        \rx_byte_cntr[2]_net_1\, C => \rx_byte_cntr[3]_net_1\, D
         => un56_sm_advance_i_cry_2_S, FCI => 
        \un58_sm_advance_i_0_data_tmp[0]\, S => OPEN, Y => OPEN, 
        FCO => \un58_sm_advance_i_0_data_tmp[1]\);
    
    RX_InProcess : SLE
      port map(D => N_311, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_InProcess\);
    
    hold_collision : SLE
      port map(D => VCC_net_1, CLK => un1_tx_collision_detect, EN
         => VCC_net_1, ALn => \N_447_i_i\, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \hold_collision\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_3\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[3]_net_1\, B => 
        un65_sm_advance_i_cry_2_S, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_2, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_3);
    
    \ReadFIFO_WR_SM.consumer_type_12[5]\ : CFG4
      generic map(INIT => x"F088")

      port map(A => RX_FIFO_DIN(3), B => N_97, C => 
        \consumer_type[5]_net_1\, D => 
        \ReadFIFO_WR_STATE[8]_net_1\, Y => \consumer_type_12[5]\);
    
    \rx_fifo_din_d1[1]\ : SLE
      port map(D => RX_FIFO_DIN(1), CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_236_i, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_fifo_din_d1[1]_net_1\);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE_3\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type4_reg(1), B => 
        consumer_type4_reg(0), C => \consumer_type[1]_net_1\, D
         => \consumer_type[0]_net_1\, Y => un38_sm_advance_i_NE_3);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE_0\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type2_reg(8), B => 
        consumer_type2_reg(7), C => \consumer_type[8]_net_1\, D
         => \consumer_type[7]_net_1\, Y => un32_sm_advance_i_NE_0);
    
    \rx_fifo_din_d3[5]\ : SLE
      port map(D => \rx_fifo_din_d2[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_236_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[5]\);
    
    rx_crc_reset : CFG2
      generic map(INIT => x"1")

      port map(A => \rx_end_rst\, B => N_480, Y => \rx_crc_reset\);
    
    \rx_fifo_din_d2[2]\ : SLE
      port map(D => \rx_fifo_din_d1[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_236_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_fifo_din_d2[2]_net_1\);
    
    \rx_byte_cntr[0]\ : SLE
      port map(D => \rx_byte_cntr_s[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_334_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_byte_cntr[0]_net_1\);
    
    \bit_cntr_RNO[2]\ : CFG4
      generic map(INIT => x"78F0")

      port map(A => \bit_cntr[0]_net_1\, B => N_265, C => 
        \bit_cntr[2]_net_1\, D => \bit_cntr[1]_net_1\, Y => 
        N_350_i_i);
    
    \rx_packet_length[0]\ : SLE
      port map(D => N_336_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_ReadFIFO_WR_STATE_14_0_0\, ALn => N_480_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_packet_length[0]_net_1\);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE_3\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type1_reg(1), B => 
        consumer_type1_reg(0), C => \consumer_type[1]_net_1\, D
         => \consumer_type[0]_net_1\, Y => un29_sm_advance_i_NE_3);
    
    \un1_rx_fifo_din_d3[2]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[2]\, B => 
        rx_crc_HighByte_en_net_1, Y => 
        \un1_rx_fifo_din_d3[2]_net_1\);
    
    \rx_packet_length_13[4]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => N_282, B => N_273, C => 
        \rx_packet_length[4]_net_1\, D => RX_FIFO_DIN(4), Y => 
        \rx_packet_length_13[4]_net_1\);
    
    \rx_crc_data_store[11]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_344_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_store[11]_net_1\);
    
    \ReadFIFO_WR_SM.consumer_type_12[2]\ : CFG4
      generic map(INIT => x"F088")

      port map(A => RX_FIFO_DIN(0), B => N_97, C => 
        \consumer_type[2]_net_1\, D => 
        \ReadFIFO_WR_STATE[8]_net_1\, Y => \consumer_type_12[2]\);
    
    \ReadFIFO_WR_STATE_ns_0_a2_0_0[6]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \hold_collision\, B => 
        \ReadFIFO_WR_STATE[5]_net_1\, C => N_236_i, Y => 
        \ReadFIFO_WR_STATE_ns_0_a2_0_0[6]_net_1\);
    
    \bit_cntr_RNO[1]\ : CFG3
      generic map(INIT => x"78")

      port map(A => \bit_cntr[0]_net_1\, B => N_265, C => 
        \bit_cntr[1]_net_1\, Y => N_326_i_i);
    
    \ReadFIFO_WR_SM.consumer_type_12[1]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => RX_FIFO_DIN(7), B => \consumer_type[1]_net_1\, 
        C => consumer_type_12_sn_N_2, D => N_670, Y => 
        \consumer_type_12[1]\);
    
    un1_ReadFIFO_WR_STATE_15_0_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => \ReadFIFO_WR_STATE[6]_net_1\, B => 
        \ReadFIFO_WR_STATE[7]_net_1\, Y => N_282);
    
    rx_end_rst_RNO : CFG2
      generic map(INIT => x"4")

      port map(A => N_582, B => idle_line, Y => N_244_i);
    
    \ReadFIFO_WR_STATE_RNI2EAL[8]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_236_i, B => \ReadFIFO_WR_STATE[8]_net_1\, Y
         => N_670);
    
    \ReadFIFO_WR_SM.consumer_type_12[7]\ : CFG4
      generic map(INIT => x"F088")

      port map(A => RX_FIFO_DIN(5), B => N_97, C => 
        \consumer_type[7]_net_1\, D => 
        \ReadFIFO_WR_STATE[8]_net_1\, Y => \consumer_type_12[7]\);
    
    \rx_crc_data_store[10]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_344_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_store[10]_net_1\);
    
    \ReadFIFO_WR_STATE_ns_i_0_a2_3_0[5]\ : CFG4
      generic map(INIT => x"010F")

      port map(A => \hold_collision\, B => 
        \ReadFIFO_WR_STATE[7]_net_1\, C => 
        \ReadFIFO_WR_STATE[4]_net_1\, D => N_236_i, Y => 
        \ReadFIFO_WR_STATE_ns_i_0_a2_3_0[5]_net_1\);
    
    \rx_byte_cntr[10]\ : SLE
      port map(D => \rx_byte_cntr_s[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_334_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_byte_cntr[10]_net_1\);
    
    un65_sm_advance_i_cry_9 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[10]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un65_sm_advance_i_cry_8\, S => un65_sm_advance_i_cry_9_S, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_9\);
    
    \SM_advancebit_cntr_RNO[2]\ : CFG4
      generic map(INIT => x"78F0")

      port map(A => \SM_advancebit_cntr[0]_net_1\, B => N_265, C
         => \SM_advancebit_cntr[2]_net_1\, D => 
        \SM_advancebit_cntr[1]_net_1\, Y => N_348_i_i);
    
    \rx_crc_data_store[7]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_330_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_store[7]_net_1\);
    
    un1_iRX_EarlyTerm_1_sqmuxa_1_0_0_a2_0 : CFG2
      generic map(INIT => x"2")

      port map(A => N_269, B => \ReadFIFO_WR_STATE[2]_net_1\, Y
         => \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0_a2_0\);
    
    \ReadFIFO_WR_SM.consumer_type_12[3]\ : CFG4
      generic map(INIT => x"F088")

      port map(A => RX_FIFO_DIN(1), B => N_97, C => 
        \consumer_type[3]_net_1\, D => 
        \ReadFIFO_WR_STATE[8]_net_1\, Y => \consumer_type_12[3]\);
    
    un56_sm_advance_i_cry_5 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[6]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un56_sm_advance_i_cry_4\, S => un56_sm_advance_i_cry_5_S, 
        Y => OPEN, FCO => \un56_sm_advance_i_cry_5\);
    
    \rx_fifo_din_d1[7]\ : SLE
      port map(D => RX_FIFO_DIN(7), CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_236_i, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_fifo_din_d1[7]_net_1\);
    
    \ReadFIFO_WR_STATE_RNO_0[4]\ : CFG4
      generic map(INIT => x"0F04")

      port map(A => \ReadFIFO_WR_STATE[9]_net_1\, B => idle_line, 
        C => \ReadFIFO_WR_STATE[8]_net_1\, D => 
        \ReadFIFO_WR_STATE_ns_i_0_a2_0_0[5]_net_1\, Y => 
        N_225_i_1);
    
    \CoreAPB3_0_APBmslave0_PREADY_i_m_i\ : CFG2
      generic map(INIT => x"D")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        CoreAPB3_0_APBmslave0_PREADY, Y => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i);
    
    \rx_byte_cntr[6]\ : SLE
      port map(D => \rx_byte_cntr_s[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_334_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_byte_cntr[6]_net_1\);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_1\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type3_reg(6), B => 
        consumer_type3_reg(5), C => \consumer_type[6]_net_1\, D
         => \consumer_type[5]_net_1\, Y => un35_sm_advance_i_NE_1);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_39\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[13]_net_1\, B => 
        \rx_crc_data_calc[12]\, C => \rx_crc_data_calc[13]\, D
         => \rx_crc_data_store[12]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[5]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[6]\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_10\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[10]_net_1\, B => 
        un65_sm_advance_i_cry_9_S, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_9, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_10);
    
    \ReadFIFO_WR_STATE[3]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \ReadFIFO_WR_STATE[3]_net_1\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_5\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[5]_net_1\, B => 
        un65_sm_advance_i_cry_4_S, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_4, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_5);
    
    \ReadFIFO_WR_STATE[1]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \ReadFIFO_WR_STATE[1]_net_1\);
    
    un56_sm_advance_i_cry_7 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[8]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un56_sm_advance_i_cry_6\, S => un56_sm_advance_i_cry_7_S, 
        Y => OPEN, FCO => \un56_sm_advance_i_cry_7\);
    
    \ReadFIFO_WR_STATE_RNI3CB2[1]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \ReadFIFO_WR_STATE[2]_net_1\, B => 
        \ReadFIFO_WR_STATE[1]_net_1\, Y => N_581);
    
    \ReadFIFO_WR_STATE[8]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \ReadFIFO_WR_STATE[8]_net_1\);
    
    \rx_crc_data_store[9]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_344_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_store[9]_net_1\);
    
    un65_sm_advance_i_cry_4 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[5]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un65_sm_advance_i_cry_3\, S => un65_sm_advance_i_cry_4_S, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_4\);
    
    \rx_byte_cntr_RNO[11]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \rx_byte_cntr[11]_net_1\, C
         => \ReadFIFO_WR_STATE_RNIHSM21_Y[9]\, D => GND_net_1, 
        FCI => \rx_byte_cntr_cry[10]\, S => \rx_byte_cntr_s[11]\, 
        Y => OPEN, FCO => OPEN);
    
    \un1_rx_fifo_din_d3[6]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[6]\, B => 
        rx_crc_HighByte_en_net_1, Y => 
        \un1_rx_fifo_din_d3[6]_net_1\);
    
    \rx_crc_data_store[4]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_330_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_store[4]_net_1\);
    
    \rx_byte_cntr[5]\ : SLE
      port map(D => \rx_byte_cntr_s[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_334_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_byte_cntr[5]_net_1\);
    
    \ReadFIFO_WR_STATE_ns_0_0[4]\ : CFG4
      generic map(INIT => x"44F0")

      port map(A => \hold_collision\, B => 
        \ReadFIFO_WR_STATE[6]_net_1\, C => 
        \ReadFIFO_WR_STATE[5]_net_1\, D => N_236_i, Y => 
        \ReadFIFO_WR_STATE_ns_0_0[4]_net_1\);
    
    \rx_fifo_din_d2[7]\ : SLE
      port map(D => \rx_fifo_din_d1[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_236_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_fifo_din_d2[7]_net_1\);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_3\ : CFG2
      generic map(INIT => x"6")

      port map(A => \consumer_type[3]_net_1\, B => 
        consumer_type4_reg(3), Y => un38_sm_advance_i_3);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_3\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type3_reg(1), B => 
        consumer_type3_reg(0), C => \consumer_type[1]_net_1\, D
         => \consumer_type[0]_net_1\, Y => un35_sm_advance_i_NE_3);
    
    \un1_rx_fifo_din_d3[3]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[3]\, B => 
        rx_crc_HighByte_en_net_1, Y => 
        \un1_rx_fifo_din_d3[3]_net_1\);
    
    \ReadFIFO_WR_STATE_RNIUBH3[3]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \ReadFIFO_WR_STATE[6]_net_1\, B => 
        \ReadFIFO_WR_STATE[5]_net_1\, C => 
        \ReadFIFO_WR_STATE[3]_net_1\, Y => 
        rx_byte_cntrlde_i_a2_0_0);
    
    \ReadFIFO_WR_STATE_ns_0[2]\ : CFG4
      generic map(INIT => x"50CC")

      port map(A => \hold_collision\, B => 
        \ReadFIFO_WR_STATE[7]_net_1\, C => 
        \ReadFIFO_WR_STATE[8]_net_1\, D => N_236_i, Y => 
        \ReadFIFO_WR_STATE_ns[2]\);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE_4\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type2_reg(9), B => 
        consumer_type2_reg(2), C => \consumer_type[9]_net_1\, D
         => \consumer_type[2]_net_1\, Y => un32_sm_advance_i_NE_4);
    
    rx_crc_LowByte_en_RNI81M61 : CFG3
      generic map(INIT => x"C8")

      port map(A => \RX_FIFO_DIN_pipe[8]\, B => N_236_i, C => 
        rx_crc_HighByte_en_net_1, Y => N_330_i);
    
    \rx_fifo_din_d3[1]\ : SLE
      port map(D => \rx_fifo_din_d2[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_236_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[1]\);
    
    un65_sm_advance_i_cry_0 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[1]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => GND_net_1, S => 
        OPEN, Y => OPEN, FCO => \un65_sm_advance_i_cry_0\);
    
    \rx_crc_data_store[2]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_330_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_store[2]_net_1\);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE_1\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type1_reg(6), B => 
        consumer_type1_reg(5), C => \consumer_type[6]_net_1\, D
         => \consumer_type[5]_net_1\, Y => un29_sm_advance_i_NE_1);
    
    \rx_packet_length_RNO[2]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => N_282, B => N_273, C => 
        \rx_packet_length[2]_net_1\, D => RX_FIFO_DIN(2), Y => 
        N_119_i);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_2\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[2]_net_1\, B => 
        un65_sm_advance_i_cry_1_S, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_1, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_2);
    
    \rx_packet_length[4]\ : SLE
      port map(D => \rx_packet_length_13[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \un1_ReadFIFO_WR_STATE_14_0_0\, 
        ALn => N_480_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[4]_net_1\);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_7\ : CFG2
      generic map(INIT => x"6")

      port map(A => \consumer_type[7]_net_1\, B => 
        consumer_type1_reg(7), Y => un29_sm_advance_i_7);
    
    N_199_i_i_o2 : CFG2
      generic map(INIT => x"8")

      port map(A => sampler_clk1x_en, B => packet_avail, Y => 
        N_265);
    
    rx_CRC_error_0_sqmuxa_0_213_a2 : CFG2
      generic map(INIT => x"8")

      port map(A => \un1_sampler_clk1x_en_0_data_tmp[7]\, B => 
        \ReadFIFO_WR_STATE[1]_net_1\, Y => N_589);
    
    un65_sm_advance_i_cry_5 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[6]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un65_sm_advance_i_cry_4\, S => un65_sm_advance_i_cry_5_S, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_5\);
    
    \rx_packet_length[1]\ : SLE
      port map(D => N_117_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_ReadFIFO_WR_STATE_14_0_0\, ALn => N_480_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_packet_length[1]_net_1\);
    
    \rx_fifo_din_d2[4]\ : SLE
      port map(D => \rx_fifo_din_d1[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_236_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_fifo_din_d2[4]_net_1\);
    
    rx_crc_reset_RNI34TD : CLKINT
      port map(A => \rx_crc_reset\, Y => rx_crc_reset_i);
    
    \rx_fifo_din_d2[3]\ : SLE
      port map(D => \rx_fifo_din_d1[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_236_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_fifo_din_d2[3]_net_1\);
    
    un65_sm_advance_i_cry_7 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[8]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un65_sm_advance_i_cry_6\, S => un65_sm_advance_i_cry_7_S, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_7\);
    
    \consumer_type[5]\ : SLE
      port map(D => \consumer_type_12[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_333_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type[5]_net_1\);
    
    \rx_crc_data_store[14]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_344_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_store[14]_net_1\);
    
    \ReadFIFO_WR_SM.consumer_type_12[8]\ : CFG4
      generic map(INIT => x"F088")

      port map(A => RX_FIFO_DIN(6), B => N_97, C => 
        \consumer_type[8]_net_1\, D => 
        \ReadFIFO_WR_STATE[8]_net_1\, Y => \consumer_type_12[8]\);
    
    \ReadFIFO_WR_SM.un40_sm_advance_i_2\ : CFG4
      generic map(INIT => x"5400")

      port map(A => DRVR_EN_c, B => un32_sm_advance_i_NE_7, C => 
        un32_sm_advance_i_NE_6, D => un30_sm_advance_i, Y => 
        un40_sm_advance_i_2);
    
    \un1_rx_fifo_din_d3[5]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[5]\, B => 
        rx_crc_HighByte_en_net_1, Y => 
        \un1_rx_fifo_din_d3[5]_net_1\);
    
    \ReadFIFO_WR_STATE[9]\ : SLE
      port map(D => N_219_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => N_480_i, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_WR_STATE[9]_net_1\);
    
    \ReadFIFO_WRITE_PROC.un15_rst_0\ : CFG3
      generic map(INIT => x"EF")

      port map(A => \RX_EarlyTerm\, B => N_480, C => clk1x_enable, 
        Y => un8_rst);
    
    \rx_byte_cntr[4]\ : SLE
      port map(D => \rx_byte_cntr_s[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_334_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_byte_cntr[4]_net_1\);
    
    \SM_advancebit_cntr[2]\ : SLE
      port map(D => N_348_i_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un8_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SM_advancebit_cntr[2]_net_1\);
    
    irx_packet_end_RNO : CFG2
      generic map(INIT => x"D")

      port map(A => N_581, B => \ReadFIFO_WR_STATE[0]_net_1\, Y
         => N_577_i);
    
    un1_ReadFIFO_WR_STATE_14_0_0_o2 : CFG2
      generic map(INIT => x"B")

      port map(A => sampler_clk1x_en, B => 
        \ReadFIFO_WR_STATE[1]_net_1\, Y => N_269);
    
    \consumer_type[0]\ : SLE
      port map(D => \consumer_type_12[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_333_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type[0]_net_1\);
    
    RX_CRC_GEN_INST : CRC16_Generator_1
      port map(RX_FIFO_DIN(7) => RX_FIFO_DIN(7), RX_FIFO_DIN(6)
         => RX_FIFO_DIN(6), RX_FIFO_DIN(5) => RX_FIFO_DIN(5), 
        RX_FIFO_DIN(4) => RX_FIFO_DIN(4), RX_FIFO_DIN(3) => 
        RX_FIFO_DIN(3), RX_FIFO_DIN(2) => RX_FIFO_DIN(2), 
        RX_FIFO_DIN(1) => RX_FIFO_DIN(1), RX_FIFO_DIN(0) => 
        RX_FIFO_DIN(0), rx_crc_data_calc(15) => 
        \rx_crc_data_calc[15]\, rx_crc_data_calc(14) => 
        \rx_crc_data_calc[14]\, rx_crc_data_calc(13) => 
        \rx_crc_data_calc[13]\, rx_crc_data_calc(12) => 
        \rx_crc_data_calc[12]\, rx_crc_data_calc(11) => 
        \rx_crc_data_calc[11]\, rx_crc_data_calc(10) => 
        \rx_crc_data_calc[10]\, rx_crc_data_calc(9) => 
        \rx_crc_data_calc[9]\, rx_crc_data_calc(8) => 
        \rx_crc_data_calc[8]\, rx_crc_data_calc(7) => 
        \rx_crc_data_calc[7]\, rx_crc_data_calc(6) => 
        \rx_crc_data_calc[6]\, rx_crc_data_calc(5) => 
        \rx_crc_data_calc[5]\, rx_crc_data_calc(4) => 
        \rx_crc_data_calc[4]\, rx_crc_data_calc(3) => 
        \rx_crc_data_calc[3]\, rx_crc_data_calc(2) => 
        \rx_crc_data_calc[2]\, rx_crc_data_calc(1) => 
        \rx_crc_data_calc[1]\, rx_crc_data_calc(0) => 
        \rx_crc_data_calc[0]\, rx_crc_gen => \rx_crc_gen\, 
        sampler_clk1x_en => sampler_clk1x_en, iRX_FIFO_wr_en => 
        iRX_FIFO_wr_en_net_1, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, rx_crc_reset_i => rx_crc_reset_i);
    
    \ReadFIFO_WR_STATE_ns_0[9]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => \ReadFIFO_WR_STATE[0]_net_1\, B => 
        \ReadFIFO_WR_STATE[1]_net_1\, C => idle_line, D => 
        sampler_clk1x_en, Y => \ReadFIFO_WR_STATE_ns[9]\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_0\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[0]_net_1\, B => 
        \rx_packet_length[0]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => GND_net_1, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_0);
    
    \ReadFIFO_WRITE_PROC.un15_rst\ : CFG2
      generic map(INIT => x"1")

      port map(A => un8_rst, B => \irx_packet_end\, Y => 
        un15_rst_i);
    
    \rx_fifo_din_d3[7]\ : SLE
      port map(D => \rx_fifo_din_d2[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_236_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[7]\);
    
    un56_sm_advance_i_cry_2 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[3]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un56_sm_advance_i_cry_1\, S => un56_sm_advance_i_cry_2_S, 
        Y => OPEN, FCO => \un56_sm_advance_i_cry_2\);
    
    \rx_packet_length[9]\ : SLE
      port map(D => N_123_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_ReadFIFO_WR_STATE_14_0_0\, ALn => N_480_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_packet_length[9]_net_1\);
    
    \rx_byte_cntr_RNI70CL6[3]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \rx_byte_cntr[3]_net_1\, C
         => \ReadFIFO_WR_STATE_RNIHSM21_Y[9]\, D => GND_net_1, 
        FCI => \rx_byte_cntr_cry[2]\, S => \rx_byte_cntr_s[3]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[3]\);
    
    \rx_fifo_din_d3[6]\ : SLE
      port map(D => \rx_fifo_din_d2[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_236_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[6]\);
    
    \rx_byte_cntr_RNIDK18C[7]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \rx_byte_cntr[7]_net_1\, C
         => \ReadFIFO_WR_STATE_RNIHSM21_Y[9]\, D => GND_net_1, 
        FCI => \rx_byte_cntr_cry[6]\, S => \rx_byte_cntr_s[7]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[7]\);
    
    rx_crc_HighByte_en_RNIG0JS : CFG2
      generic map(INIT => x"8")

      port map(A => N_236_i, B => rx_crc_HighByte_en_net_1, Y => 
        N_344_i);
    
    \consumer_type[9]\ : SLE
      port map(D => \consumer_type_12[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_333_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type[9]_net_1\);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_6\ : CFG4
      generic map(INIT => x"FFF6")

      port map(A => \consumer_type[4]_net_1\, B => 
        consumer_type3_reg(4), C => un35_sm_advance_i_NE_3, D => 
        un35_sm_advance_i_3, Y => un35_sm_advance_i_NE_6);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_33\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[11]_net_1\, B => 
        \rx_crc_data_calc[10]\, C => \rx_crc_data_calc[11]\, D
         => \rx_crc_data_store[10]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[4]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[5]\);
    
    \rx_crc_data_store[6]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_330_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_store[6]_net_1\);
    
    ReadFIFO_WR_STATE_1_sqmuxa_1_0_a3_0_a2 : CFG3
      generic map(INIT => x"04")

      port map(A => \hold_collision\, B => 
        \ReadFIFO_WR_STATE[5]_net_1\, C => 
        \un58_sm_advance_i_0_data_tmp[5]\, Y => 
        ReadFIFO_WR_STATE_1_sqmuxa_1);
    
    SM_advance_i_RNIAH4K : CFG2
      generic map(INIT => x"8")

      port map(A => sampler_clk1x_en, B => \SM_advance_i\, Y => 
        N_236_i);
    
    \ReadFIFO_WR_STATE_ns_0[4]\ : CFG4
      generic map(INIT => x"F4F0")

      port map(A => \hold_collision\, B => 
        \ReadFIFO_WR_STATE[5]_net_1\, C => 
        \ReadFIFO_WR_STATE_ns_0_0[4]_net_1\, D => 
        \un58_sm_advance_i_0_data_tmp[5]\, Y => 
        \ReadFIFO_WR_STATE_ns[4]\);
    
    SM_advance_i : SLE
      port map(D => un2_packet_avail, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_265, ALn => un8_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SM_advance_i\);
    
    \ReadFIFO_WR_STATE_ns_0[1]\ : CFG3
      generic map(INIT => x"DC")

      port map(A => N_236_i, B => N_396, C => 
        \ReadFIFO_WR_STATE[8]_net_1\, Y => 
        \ReadFIFO_WR_STATE_ns[1]\);
    
    un65_sm_advance_i_cry_8 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \rx_packet_length[9]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un65_sm_advance_i_cry_7\, S => un65_sm_advance_i_cry_8_S, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_8\);
    
    \consumer_type[3]\ : SLE
      port map(D => \consumer_type_12[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_333_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type[3]_net_1\);
    
    \rx_byte_cntr[3]\ : SLE
      port map(D => \rx_byte_cntr_s[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_334_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_byte_cntr[3]_net_1\);
    
    RX_InProcess_d1_RNIKPES : CFG3
      generic map(INIT => x"80")

      port map(A => RX_InProcess_d1_net_1, B => 
        iRX_FIFO_wr_en_net_1, C => sampler_clk1x_en, Y => N_366_i);
    
    \rx_crc_data_store[3]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_330_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_store[3]_net_1\);
    
    \rx_byte_cntr[7]\ : SLE
      port map(D => \rx_byte_cntr_s[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_334_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_byte_cntr[7]_net_1\);
    
    \RX_InProcess_d1\ : SLE
      port map(D => \RX_InProcess\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        RX_InProcess_d1_net_1);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE_5\ : CFG4
      generic map(INIT => x"FFF6")

      port map(A => \consumer_type[8]_net_1\, B => 
        consumer_type1_reg(8), C => un29_sm_advance_i_NE_1, D => 
        un29_sm_advance_i_7, Y => un29_sm_advance_i_NE_5);
    
    \consumer_type[8]\ : SLE
      port map(D => \consumer_type_12[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_333_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type[8]_net_1\);
    
    \rx_packet_length[3]\ : SLE
      port map(D => \rx_packet_length_13[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \un1_ReadFIFO_WR_STATE_14_0_0\, 
        ALn => N_480_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[3]_net_1\);
    
    \SM_advancebit_cntr_RNO[1]\ : CFG3
      generic map(INIT => x"78")

      port map(A => \SM_advancebit_cntr[0]_net_1\, B => N_265, C
         => \SM_advancebit_cntr[1]_net_1\, Y => N_325_i_i);
    
    irx_packet_end : SLE
      port map(D => N_577_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \irx_packet_end\);
    
    rx_crc_gen : SLE
      port map(D => un1_ReadFIFO_WR_STATE_15, CLK => 
        CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_gen\);
    
    \rx_byte_cntr_RNIMKC1F[9]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \rx_byte_cntr[9]_net_1\, C
         => \ReadFIFO_WR_STATE_RNIHSM21_Y[9]\, D => GND_net_1, 
        FCI => \rx_byte_cntr_cry[8]\, S => \rx_byte_cntr_s[9]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[9]\);
    
    \ReadFIFO_WRITE_PROC.un15_rst_0_RNIR373\ : CFG1
      generic map(INIT => "01")

      port map(A => un8_rst, Y => un8_rst_i);
    
    \rx_fifo_din_d1[6]\ : SLE
      port map(D => RX_FIFO_DIN(6), CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_236_i, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_fifo_din_d1[6]_net_1\);
    
    \rx_packet_length_13[7]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => N_282, B => N_273, C => 
        \rx_packet_length[7]_net_1\, D => RX_FIFO_DIN(7), Y => 
        \rx_packet_length_13[7]_net_1\);
    
    \rx_fifo_din_d3[3]\ : SLE
      port map(D => \rx_fifo_din_d2[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_236_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[3]\);
    
    un1_ReadFIFO_WR_STATE_14_0_0_a2 : CFG4
      generic map(INIT => x"1000")

      port map(A => \ReadFIFO_WR_STATE[3]_net_1\, B => 
        \ReadFIFO_WR_STATE[5]_net_1\, C => N_269, D => 
        un1_ReadFIFO_WR_STATE_14_0_0_a2_0, Y => N_405);
    
    \rx_fifo_din_d3[0]\ : SLE
      port map(D => \rx_fifo_din_d2[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_236_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[0]\);
    
    \ReadFIFO_WR_STATE[5]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \ReadFIFO_WR_STATE[5]_net_1\);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_1\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[1]_net_1\, B => 
        \rx_crc_data_calc[0]\, C => \rx_crc_data_calc[1]\, D => 
        \rx_crc_data_store[0]_net_1\, FCI => GND_net_1, S => OPEN, 
        Y => OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[0]\);
    
    un65_sm_advance_i_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_packet_length[2]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \un65_sm_advance_i_cry_0\, S => un65_sm_advance_i_cry_1_S, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_1\);
    
    rx_packet_complt_RNIF8T4 : CFG1
      generic map(INIT => "01")

      port map(A => rx_packet_complt_net_1, Y => 
        rx_packet_complt_i);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_3\ : CFG2
      generic map(INIT => x"6")

      port map(A => \consumer_type[3]_net_1\, B => 
        consumer_type2_reg(3), Y => un32_sm_advance_i_3);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_27\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[7]_net_1\, B => 
        \rx_crc_data_calc[6]\, C => \rx_crc_data_calc[7]\, D => 
        \rx_crc_data_store[6]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[2]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[3]\);
    
    \consumer_type[2]\ : SLE
      port map(D => \consumer_type_12[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_333_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type[2]_net_1\);
    
    \ReadFIFO_WR_STATE_ns_0[7]\ : CFG4
      generic map(INIT => x"50CC")

      port map(A => \hold_collision\, B => 
        \ReadFIFO_WR_STATE[2]_net_1\, C => 
        \ReadFIFO_WR_STATE[3]_net_1\, D => N_236_i, Y => 
        \ReadFIFO_WR_STATE_ns[7]\);
    
    \rx_byte_cntr_RNINB128[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \rx_byte_cntr[4]_net_1\, C
         => \ReadFIFO_WR_STATE_RNIHSM21_Y[9]\, D => GND_net_1, 
        FCI => \rx_byte_cntr_cry[3]\, S => \rx_byte_cntr_s[4]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[4]\);
    
    \rx_crc_data_store[15]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_344_i, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_store[15]_net_1\);
    
    rx_CRC_error_RNIASV4 : CFG1
      generic map(INIT => "01")

      port map(A => rx_CRC_error_net_1, Y => rx_CRC_error_i);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE_3\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type2_reg(1), B => 
        consumer_type2_reg(0), C => \consumer_type[1]_net_1\, D
         => \consumer_type[0]_net_1\, Y => un32_sm_advance_i_NE_3);
    
    \rx_packet_length_RNO[0]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => N_282, B => N_273, C => 
        \rx_packet_length[0]_net_1\, D => RX_FIFO_DIN(0), Y => 
        N_336_i);
    
    rx_end_rst_0_sqmuxa_i_o3_0_a2 : CFG2
      generic map(INIT => x"1")

      port map(A => \ReadFIFO_WR_STATE[4]_net_1\, B => 
        \ReadFIFO_WR_STATE[0]_net_1\, Y => N_582);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity AFE_RX_SM is

    port( RX_FIFO_DIN          : in    std_logic_vector(7 downto 0);
          manches_in_dly       : in    std_logic_vector(1 downto 0);
          irx_center_sample    : in    std_logic;
          RX_EarlyTerm         : in    std_logic;
          N_480                : in    std_logic;
          idle_line            : in    std_logic;
          long_reset           : in    std_logic;
          CommsFPGA_CCC_0_LOCK : in    std_logic;
          clk1x_enable         : out   std_logic;
          packet_avail         : out   std_logic;
          N_480_i              : in    std_logic;
          CommsFPGA_CCC_0_GL0  : in    std_logic;
          N_584_i_i            : out   std_logic
        );

end AFE_RX_SM;

architecture DEF_ARCH of AFE_RX_SM is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_584_i, \irx_packet_end_all_RNIB6KE\, 
        \start_bit_mask\, VCC_net_1, \start_bit_mask_1\, 
        \start_bit_maskce\, GND_net_1, \RX_EarlyTerm_s\, 
        \RX_EarlyTerm_s_0\, \start_bit_cntr[0]_net_1\, N_12_i, 
        \start_bit_cntr[1]_net_1\, N_10_i, 
        \start_bit_cntr[2]_net_1\, N_8_i, 
        \start_bit_cntr[3]_net_1\, N_6_i, \AFE_RX_STATE[4]_net_1\, 
        N_76_i, \AFE_RX_STATE[3]_net_1\, \AFE_RX_STATE_ns[1]\, 
        \AFE_RX_STATE[2]_net_1\, \AFE_RX_STATE_ns[2]_net_1\, 
        \packet_avail\, \AFE_RX_STATE_11[1]\, 
        \AFE_RX_STATE[0]_net_1\, \AFE_RX_STATE_ns[4]\, 
        rx_packet_end_all, irx_packet_end_all_4, clk1x_enable_6, 
        N_356, clk1x_enable_6_0_0_1, 
        \AFE_RX_STATE_ns_a4_0_a2_0_2[3]_net_1\, 
        \AFE_RX_STATE_ns_a4_0_a2_0_1[3]\, N_392_6, N_280, N_367, 
        \start_bit_cntr_0_i_0_0[1]_net_1\, N_392, un1_rx_fifo_din
         : std_logic;

begin 

    packet_avail <= \packet_avail\;

    \AFE_RX_STATE_ns_i_0_a2_0[0]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \AFE_RX_STATE[4]_net_1\, B => 
        manches_in_dly(0), C => manches_in_dly(1), Y => 
        \AFE_RX_STATE_ns[1]\);
    
    \start_bit_cntr[2]\ : SLE
      port map(D => N_8_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[2]_net_1\);
    
    RX_EarlyTerm_s_0 : CFG2
      generic map(INIT => x"4")

      port map(A => N_480, B => RX_EarlyTerm, Y => 
        \RX_EarlyTerm_s_0\);
    
    \AFE_RX_STATE[3]\ : SLE
      port map(D => \AFE_RX_STATE_ns[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \AFE_RX_STATE[3]_net_1\);
    
    irx_packet_end_all_RNIB6KE : CFG3
      generic map(INIT => x"FB")

      port map(A => rx_packet_end_all, B => CommsFPGA_CCC_0_LOCK, 
        C => long_reset, Y => \irx_packet_end_all_RNIB6KE\);
    
    irx_packet_end_all_RNIB6KE_0 : CLKINT
      port map(A => \irx_packet_end_all_RNIB6KE\, Y => N_584_i);
    
    \AFE_RX_SM.un1_rx_fifo_din_0_a2_1\ : CFG3
      generic map(INIT => x"10")

      port map(A => RX_FIFO_DIN(3), B => RX_FIFO_DIN(2), C => 
        RX_FIFO_DIN(0), Y => \AFE_RX_STATE_ns_a4_0_a2_0_1[3]\);
    
    irx_packet_end_all_RNIB6KE_1 : CFG1
      generic map(INIT => "01")

      port map(A => N_584_i, Y => N_584_i_i);
    
    \start_bit_cntr_0_i_0_0[1]\ : CFG4
      generic map(INIT => x"CDCF")

      port map(A => irx_center_sample, B => N_584_i, C => 
        \start_bit_cntr[1]_net_1\, D => \start_bit_cntr[0]_net_1\, 
        Y => \start_bit_cntr_0_i_0_0[1]_net_1\);
    
    \AFE_RX_STATE_ns[2]\ : CFG4
      generic map(INIT => x"5150")

      port map(A => idle_line, B => un1_rx_fifo_din, C => 
        \AFE_RX_STATE[3]_net_1\, D => \AFE_RX_STATE[2]_net_1\, Y
         => \AFE_RX_STATE_ns[2]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \start_bit_cntr_0_i_0_o2[0]\ : CFG3
      generic map(INIT => x"FB")

      port map(A => \start_bit_cntr[2]_net_1\, B => 
        \start_bit_cntr[1]_net_1\, C => \start_bit_cntr[3]_net_1\, 
        Y => N_367);
    
    start_bit_maskce : CFG4
      generic map(INIT => x"FFFE")

      port map(A => N_480, B => N_584_i, C => rx_packet_end_all, 
        D => irx_center_sample, Y => \start_bit_maskce\);
    
    \start_bit_cntr[3]\ : SLE
      port map(D => N_6_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[3]_net_1\);
    
    \start_bit_cntr_RNO[3]\ : CFG4
      generic map(INIT => x"2130")

      port map(A => N_280, B => N_584_i, C => 
        \start_bit_cntr[3]_net_1\, D => \start_bit_cntr[2]_net_1\, 
        Y => N_6_i);
    
    \AFE_RX_STATE_ns_a4_0[3]\ : CFG4
      generic map(INIT => x"FF04")

      port map(A => \RX_EarlyTerm_s\, B => \packet_avail\, C => 
        idle_line, D => N_392, Y => \AFE_RX_STATE_11[1]\);
    
    \AFE_RX_STATE[1]\ : SLE
      port map(D => \AFE_RX_STATE_11[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \packet_avail\);
    
    \AFE_RX_STATE[4]\ : SLE
      port map(D => N_76_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => N_480_i, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \AFE_RX_STATE[4]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \start_bit_cntr[0]\ : SLE
      port map(D => N_12_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[0]_net_1\);
    
    \start_bit_cntr_RNO[2]\ : CFG4
      generic map(INIT => x"2210")

      port map(A => N_280, B => N_584_i, C => 
        \start_bit_cntr[3]_net_1\, D => \start_bit_cntr[2]_net_1\, 
        Y => N_8_i);
    
    RX_EarlyTerm_s : SLE
      port map(D => \RX_EarlyTerm_s_0\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_EarlyTerm_s\);
    
    \start_bit_cntr[1]\ : SLE
      port map(D => N_10_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[1]_net_1\);
    
    \AFE_RX_STATE_RNO[4]\ : CFG3
      generic map(INIT => x"54")

      port map(A => \AFE_RX_STATE_ns[1]\, B => 
        \AFE_RX_STATE[4]_net_1\, C => idle_line, Y => N_76_i);
    
    \AFE_RX_STATE[0]\ : SLE
      port map(D => \AFE_RX_STATE_ns[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \AFE_RX_STATE[0]_net_1\);
    
    \AFE_RX_SM.un1_rx_fifo_din_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => RX_FIFO_DIN(1), B => RX_FIFO_DIN(6), C => 
        N_392_6, D => \AFE_RX_STATE_ns_a4_0_a2_0_1[3]\, Y => 
        un1_rx_fifo_din);
    
    \AFE_RX_STATE_ns_a4_0_a2_0[3]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \AFE_RX_STATE_ns_a4_0_a2_0_2[3]_net_1\, B => 
        \AFE_RX_STATE_ns_a4_0_a2_0_1[3]\, C => N_392_6, Y => 
        N_392);
    
    \start_bit_cntr_RNO[0]\ : CFG4
      generic map(INIT => x"1330")

      port map(A => N_367, B => N_584_i, C => 
        \start_bit_cntr[0]_net_1\, D => irx_center_sample, Y => 
        N_12_i);
    
    start_bit_mask_1 : CFG4
      generic map(INIT => x"EFCC")

      port map(A => N_367, B => N_584_i, C => 
        \start_bit_cntr[0]_net_1\, D => irx_center_sample, Y => 
        \start_bit_mask_1\);
    
    \AFE_RX_SM.un1_rx_fifo_din_0_a2_5\ : CFG4
      generic map(INIT => x"0100")

      port map(A => RX_FIFO_DIN(5), B => RX_FIFO_DIN(4), C => 
        \start_bit_mask\, D => RX_FIFO_DIN(7), Y => N_392_6);
    
    \AFE_RX_STATE_ns_0[4]\ : CFG4
      generic map(INIT => x"00EC")

      port map(A => \RX_EarlyTerm_s\, B => 
        \AFE_RX_STATE[0]_net_1\, C => \packet_avail\, D => 
        idle_line, Y => \AFE_RX_STATE_ns[4]\);
    
    \AFE_RX_SM.clk1x_enable_6_0_0\ : CFG4
      generic map(INIT => x"F4FB")

      port map(A => N_356, B => clk1x_enable_6_0_0_1, C => 
        \AFE_RX_STATE[0]_net_1\, D => idle_line, Y => 
        clk1x_enable_6);
    
    \AFE_RX_SM.irx_packet_end_all_4_0_a4_0_a2\ : CFG2
      generic map(INIT => x"2")

      port map(A => idle_line, B => \AFE_RX_STATE[4]_net_1\, Y
         => irx_packet_end_all_4);
    
    \AFE_RX_SM.clk1x_enable_6_0_0_1\ : CFG4
      generic map(INIT => x"0603")

      port map(A => manches_in_dly(1), B => idle_line, C => 
        \packet_avail\, D => manches_in_dly(0), Y => 
        clk1x_enable_6_0_0_1);
    
    \start_bit_cntr_RNO[1]\ : CFG4
      generic map(INIT => x"00F1")

      port map(A => \start_bit_cntr[3]_net_1\, B => 
        \start_bit_cntr[2]_net_1\, C => N_280, D => 
        \start_bit_cntr_0_i_0_0[1]_net_1\, Y => N_10_i);
    
    \AFE_RX_STATE_ns_a4_0_a2_0_2[3]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => idle_line, B => \AFE_RX_STATE[2]_net_1\, C
         => RX_FIFO_DIN(1), D => RX_FIFO_DIN(6), Y => 
        \AFE_RX_STATE_ns_a4_0_a2_0_2[3]_net_1\);
    
    irx_packet_end_all : SLE
      port map(D => irx_packet_end_all_4, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rx_packet_end_all);
    
    \AFE_RX_SM.clk1x_enable_6_0_0_o2\ : CFG2
      generic map(INIT => x"E")

      port map(A => \AFE_RX_STATE[2]_net_1\, B => 
        \AFE_RX_STATE[3]_net_1\, Y => N_356);
    
    \AFE_RX_STATE[2]\ : SLE
      port map(D => \AFE_RX_STATE_ns[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => N_480_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \AFE_RX_STATE[2]_net_1\);
    
    start_bit_mask : SLE
      port map(D => \start_bit_mask_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \start_bit_maskce\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \start_bit_mask\);
    
    \clk1x_enable\ : SLE
      port map(D => clk1x_enable_6, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        clk1x_enable);
    
    \start_bit_cntr_0_i_0_o2_0[3]\ : CFG3
      generic map(INIT => x"7F")

      port map(A => \start_bit_cntr[0]_net_1\, B => 
        irx_center_sample, C => \start_bit_cntr[1]_net_1\, Y => 
        N_280);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity ManchesDecoder is

    port( RX_FIFO_DIN_pipe                   : out   std_logic_vector(8 downto 0);
          consumer_type1_reg                 : in    std_logic_vector(9 downto 0);
          consumer_type2_reg                 : in    std_logic_vector(9 downto 0);
          consumer_type3_reg                 : in    std_logic_vector(9 downto 0);
          consumer_type4_reg                 : in    std_logic_vector(9 downto 0);
          RX_FIFO_DIN                        : out   std_logic_vector(7 downto 0);
          manches_in_dly                     : out   std_logic_vector(1 downto 0);
          rx_CRC_error                       : out   std_logic;
          rx_CRC_error_i                     : out   std_logic;
          rx_packet_complt                   : out   std_logic;
          rx_packet_complt_i                 : out   std_logic;
          rx_crc_HighByte_en                 : out   std_logic;
          iRX_FIFO_wr_en                     : out   std_logic;
          RX_InProcess_d1                    : out   std_logic;
          TX_collision_detect                : in    std_logic;
          tx_col_detect_en                   : in    std_logic;
          CoreAPB3_0_APBmslave0_PSELx        : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY       : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY_i_m_i : out   std_logic;
          N_366_i                            : out   std_logic;
          DRVR_EN_c                          : in    std_logic;
          CommsFPGA_CCC_0_LOCK               : in    std_logic;
          long_reset                         : in    std_logic;
          N_480                              : in    std_logic;
          RX_EarlyTerm                       : out   std_logic;
          CommsFPGA_CCC_0_GL0                : in    std_logic;
          N_480_i                            : in    std_logic;
          sampler_clk1x_en                   : out   std_logic;
          MANCH_OUT_P_c                      : in    std_logic;
          MANCHESTER_IN_c                    : in    std_logic;
          internal_loopback                  : in    std_logic;
          N_268_i                            : in    std_logic
        );

end ManchesDecoder;

architecture DEF_ARCH of ManchesDecoder is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component ManchesDecoder_Adapter
    port( manches_in_dly      : out   std_logic_vector(1 downto 0);
          RX_FIFO_DIN         : out   std_logic_vector(7 downto 0);
          idle_line           : out   std_logic;
          N_268_i             : in    std_logic := 'U';
          internal_loopback   : in    std_logic := 'U';
          MANCHESTER_IN_c     : in    std_logic := 'U';
          MANCH_OUT_P_c       : in    std_logic := 'U';
          irx_center_sample   : out   std_logic;
          N_447_i_i           : in    std_logic := 'U';
          sampler_clk1x_en    : out   std_logic;
          N_480_i             : in    std_logic := 'U';
          clk1x_enable        : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          N_584_i_i           : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component ReadFIFO_Write_SM
    port( consumer_type4_reg                 : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type3_reg                 : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type2_reg                 : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type1_reg                 : in    std_logic_vector(9 downto 0) := (others => 'U');
          RX_FIFO_DIN                        : in    std_logic_vector(7 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe                   : out   std_logic_vector(8 downto 0);
          DRVR_EN_c                          : in    std_logic := 'U';
          N_366_i                            : out   std_logic;
          clk1x_enable                       : in    std_logic := 'U';
          N_480                              : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY_i_m_i : out   std_logic;
          CoreAPB3_0_APBmslave0_PREADY       : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PSELx        : in    std_logic := 'U';
          tx_col_detect_en                   : in    std_logic := 'U';
          TX_collision_detect                : in    std_logic := 'U';
          sampler_clk1x_en                   : in    std_logic := 'U';
          idle_line                          : in    std_logic := 'U';
          packet_avail                       : in    std_logic := 'U';
          N_447_i_i                          : out   std_logic;
          RX_InProcess_d1                    : out   std_logic;
          iRX_FIFO_wr_en                     : out   std_logic;
          RX_EarlyTerm                       : out   std_logic;
          rx_crc_HighByte_en                 : out   std_logic;
          CommsFPGA_CCC_0_GL0                : in    std_logic := 'U';
          N_480_i                            : in    std_logic := 'U';
          rx_packet_complt_i                 : out   std_logic;
          rx_packet_complt                   : out   std_logic;
          rx_CRC_error_i                     : out   std_logic;
          rx_CRC_error                       : out   std_logic
        );
  end component;

  component AFE_RX_SM
    port( RX_FIFO_DIN          : in    std_logic_vector(7 downto 0) := (others => 'U');
          manches_in_dly       : in    std_logic_vector(1 downto 0) := (others => 'U');
          irx_center_sample    : in    std_logic := 'U';
          RX_EarlyTerm         : in    std_logic := 'U';
          N_480                : in    std_logic := 'U';
          idle_line            : in    std_logic := 'U';
          long_reset           : in    std_logic := 'U';
          CommsFPGA_CCC_0_LOCK : in    std_logic := 'U';
          clk1x_enable         : out   std_logic;
          packet_avail         : out   std_logic;
          N_480_i              : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0  : in    std_logic := 'U';
          N_584_i_i            : out   std_logic
        );
  end component;

    signal \manches_in_dly[0]\, \manches_in_dly[1]\, 
        \RX_FIFO_DIN[0]\, \RX_FIFO_DIN[1]\, \RX_FIFO_DIN[2]\, 
        \RX_FIFO_DIN[3]\, \RX_FIFO_DIN[4]\, \RX_FIFO_DIN[5]\, 
        \RX_FIFO_DIN[6]\, \RX_FIFO_DIN[7]\, idle_line, 
        irx_center_sample, N_447_i_i, \sampler_clk1x_en\, 
        clk1x_enable, N_584_i_i, \RX_EarlyTerm\, packet_avail, 
        GND_net_1, VCC_net_1 : std_logic;

    for all : ManchesDecoder_Adapter
	Use entity work.ManchesDecoder_Adapter(DEF_ARCH);
    for all : ReadFIFO_Write_SM
	Use entity work.ReadFIFO_Write_SM(DEF_ARCH);
    for all : AFE_RX_SM
	Use entity work.AFE_RX_SM(DEF_ARCH);
begin 

    RX_FIFO_DIN(7) <= \RX_FIFO_DIN[7]\;
    RX_FIFO_DIN(6) <= \RX_FIFO_DIN[6]\;
    RX_FIFO_DIN(5) <= \RX_FIFO_DIN[5]\;
    RX_FIFO_DIN(4) <= \RX_FIFO_DIN[4]\;
    RX_FIFO_DIN(3) <= \RX_FIFO_DIN[3]\;
    RX_FIFO_DIN(2) <= \RX_FIFO_DIN[2]\;
    RX_FIFO_DIN(1) <= \RX_FIFO_DIN[1]\;
    RX_FIFO_DIN(0) <= \RX_FIFO_DIN[0]\;
    manches_in_dly(1) <= \manches_in_dly[1]\;
    manches_in_dly(0) <= \manches_in_dly[0]\;
    RX_EarlyTerm <= \RX_EarlyTerm\;
    sampler_clk1x_en <= \sampler_clk1x_en\;

    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    MANCHESTER_DECODER_ADAPTER_INST : ManchesDecoder_Adapter
      port map(manches_in_dly(1) => \manches_in_dly[1]\, 
        manches_in_dly(0) => \manches_in_dly[0]\, RX_FIFO_DIN(7)
         => \RX_FIFO_DIN[7]\, RX_FIFO_DIN(6) => \RX_FIFO_DIN[6]\, 
        RX_FIFO_DIN(5) => \RX_FIFO_DIN[5]\, RX_FIFO_DIN(4) => 
        \RX_FIFO_DIN[4]\, RX_FIFO_DIN(3) => \RX_FIFO_DIN[3]\, 
        RX_FIFO_DIN(2) => \RX_FIFO_DIN[2]\, RX_FIFO_DIN(1) => 
        \RX_FIFO_DIN[1]\, RX_FIFO_DIN(0) => \RX_FIFO_DIN[0]\, 
        idle_line => idle_line, N_268_i => N_268_i, 
        internal_loopback => internal_loopback, MANCHESTER_IN_c
         => MANCHESTER_IN_c, MANCH_OUT_P_c => MANCH_OUT_P_c, 
        irx_center_sample => irx_center_sample, N_447_i_i => 
        N_447_i_i, sampler_clk1x_en => \sampler_clk1x_en\, 
        N_480_i => N_480_i, clk1x_enable => clk1x_enable, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, N_584_i_i => 
        N_584_i_i);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    ReadFIFO_Write_SM_PROC : ReadFIFO_Write_SM
      port map(consumer_type4_reg(9) => consumer_type4_reg(9), 
        consumer_type4_reg(8) => consumer_type4_reg(8), 
        consumer_type4_reg(7) => consumer_type4_reg(7), 
        consumer_type4_reg(6) => consumer_type4_reg(6), 
        consumer_type4_reg(5) => consumer_type4_reg(5), 
        consumer_type4_reg(4) => consumer_type4_reg(4), 
        consumer_type4_reg(3) => consumer_type4_reg(3), 
        consumer_type4_reg(2) => consumer_type4_reg(2), 
        consumer_type4_reg(1) => consumer_type4_reg(1), 
        consumer_type4_reg(0) => consumer_type4_reg(0), 
        consumer_type3_reg(9) => consumer_type3_reg(9), 
        consumer_type3_reg(8) => consumer_type3_reg(8), 
        consumer_type3_reg(7) => consumer_type3_reg(7), 
        consumer_type3_reg(6) => consumer_type3_reg(6), 
        consumer_type3_reg(5) => consumer_type3_reg(5), 
        consumer_type3_reg(4) => consumer_type3_reg(4), 
        consumer_type3_reg(3) => consumer_type3_reg(3), 
        consumer_type3_reg(2) => consumer_type3_reg(2), 
        consumer_type3_reg(1) => consumer_type3_reg(1), 
        consumer_type3_reg(0) => consumer_type3_reg(0), 
        consumer_type2_reg(9) => consumer_type2_reg(9), 
        consumer_type2_reg(8) => consumer_type2_reg(8), 
        consumer_type2_reg(7) => consumer_type2_reg(7), 
        consumer_type2_reg(6) => consumer_type2_reg(6), 
        consumer_type2_reg(5) => consumer_type2_reg(5), 
        consumer_type2_reg(4) => consumer_type2_reg(4), 
        consumer_type2_reg(3) => consumer_type2_reg(3), 
        consumer_type2_reg(2) => consumer_type2_reg(2), 
        consumer_type2_reg(1) => consumer_type2_reg(1), 
        consumer_type2_reg(0) => consumer_type2_reg(0), 
        consumer_type1_reg(9) => consumer_type1_reg(9), 
        consumer_type1_reg(8) => consumer_type1_reg(8), 
        consumer_type1_reg(7) => consumer_type1_reg(7), 
        consumer_type1_reg(6) => consumer_type1_reg(6), 
        consumer_type1_reg(5) => consumer_type1_reg(5), 
        consumer_type1_reg(4) => consumer_type1_reg(4), 
        consumer_type1_reg(3) => consumer_type1_reg(3), 
        consumer_type1_reg(2) => consumer_type1_reg(2), 
        consumer_type1_reg(1) => consumer_type1_reg(1), 
        consumer_type1_reg(0) => consumer_type1_reg(0), 
        RX_FIFO_DIN(7) => \RX_FIFO_DIN[7]\, RX_FIFO_DIN(6) => 
        \RX_FIFO_DIN[6]\, RX_FIFO_DIN(5) => \RX_FIFO_DIN[5]\, 
        RX_FIFO_DIN(4) => \RX_FIFO_DIN[4]\, RX_FIFO_DIN(3) => 
        \RX_FIFO_DIN[3]\, RX_FIFO_DIN(2) => \RX_FIFO_DIN[2]\, 
        RX_FIFO_DIN(1) => \RX_FIFO_DIN[1]\, RX_FIFO_DIN(0) => 
        \RX_FIFO_DIN[0]\, RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), DRVR_EN_c => DRVR_EN_c, N_366_i => 
        N_366_i, clk1x_enable => clk1x_enable, N_480 => N_480, 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, 
        CoreAPB3_0_APBmslave0_PREADY => 
        CoreAPB3_0_APBmslave0_PREADY, CoreAPB3_0_APBmslave0_PSELx
         => CoreAPB3_0_APBmslave0_PSELx, tx_col_detect_en => 
        tx_col_detect_en, TX_collision_detect => 
        TX_collision_detect, sampler_clk1x_en => 
        \sampler_clk1x_en\, idle_line => idle_line, packet_avail
         => packet_avail, N_447_i_i => N_447_i_i, RX_InProcess_d1
         => RX_InProcess_d1, iRX_FIFO_wr_en => iRX_FIFO_wr_en, 
        RX_EarlyTerm => \RX_EarlyTerm\, rx_crc_HighByte_en => 
        rx_crc_HighByte_en, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, N_480_i => N_480_i, 
        rx_packet_complt_i => rx_packet_complt_i, 
        rx_packet_complt => rx_packet_complt, rx_CRC_error_i => 
        rx_CRC_error_i, rx_CRC_error => rx_CRC_error);
    
    AFE_RX_STATE_MACHINE : AFE_RX_SM
      port map(RX_FIFO_DIN(7) => \RX_FIFO_DIN[7]\, RX_FIFO_DIN(6)
         => \RX_FIFO_DIN[6]\, RX_FIFO_DIN(5) => \RX_FIFO_DIN[5]\, 
        RX_FIFO_DIN(4) => \RX_FIFO_DIN[4]\, RX_FIFO_DIN(3) => 
        \RX_FIFO_DIN[3]\, RX_FIFO_DIN(2) => \RX_FIFO_DIN[2]\, 
        RX_FIFO_DIN(1) => \RX_FIFO_DIN[1]\, RX_FIFO_DIN(0) => 
        \RX_FIFO_DIN[0]\, manches_in_dly(1) => 
        \manches_in_dly[1]\, manches_in_dly(0) => 
        \manches_in_dly[0]\, irx_center_sample => 
        irx_center_sample, RX_EarlyTerm => \RX_EarlyTerm\, N_480
         => N_480, idle_line => idle_line, long_reset => 
        long_reset, CommsFPGA_CCC_0_LOCK => CommsFPGA_CCC_0_LOCK, 
        clk1x_enable => clk1x_enable, packet_avail => 
        packet_avail, N_480_i => N_480_i, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, N_584_i_i => N_584_i_i);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top is

    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0);
          fifo_MEMRADDR             : in    std_logic_vector(12 downto 0);
          fifo_MEMWE                : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          N_283_i                   : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component RAM1K18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_CLK         : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ARST_N      : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          A_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_CLK         : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ARST_N      : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          B_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_WMODE       : in    std_logic := 'U';
          B_EN          : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_WMODE       : in    std_logic := 'U';
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;
    signal nc151, nc23, nc58, nc116, nc74, nc133, nc167, nc84, 
        nc39, nc72, nc82, nc145, nc160, nc57, nc156, nc125, nc73, 
        nc107, nc66, nc83, nc9, nc171, nc54, nc135, nc41, nc100, 
        nc52, nc29, nc118, nc60, nc141, nc45, nc53, nc121, nc158, 
        nc162, nc11, nc131, nc96, nc79, nc146, nc89, nc119, nc48, 
        nc126, nc15, nc102, nc3, nc47, nc90, nc159, nc136, nc59, 
        nc18, nc44, nc117, nc164, nc148, nc42, nc17, nc2, nc110, 
        nc128, nc43, nc157, nc36, nc61, nc104, nc138, nc14, nc150, 
        nc149, nc12, nc30, nc65, nc7, nc129, nc8, nc13, nc26, 
        nc139, nc163, nc112, nc68, nc49, nc170, nc91, nc5, nc20, 
        nc147, nc67, nc152, nc127, nc103, nc76, nc140, nc86, nc95, 
        nc120, nc165, nc137, nc64, nc19, nc70, nc62, nc80, nc130, 
        nc98, nc114, nc56, nc105, nc63, nc97, nc161, nc31, nc154, 
        nc50, nc142, nc94, nc122, nc35, nc4, nc92, nc101, nc166, 
        nc132, nc21, nc93, nc69, nc38, nc113, nc106, nc25, nc1, 
        nc37, nc144, nc153, nc46, nc71, nc124, nc81, nc168, nc34, 
        nc28, nc115, nc134, nc32, nc40, nc99, nc75, nc85, nc27, 
        nc108, nc16, nc155, nc51, nc33, nc169, nc78, nc24, nc88, 
        nc111, nc55, nc10, nc22, nc143, nc77, nc6, nc109, nc87, 
        nc123 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C2 : RAM1K18
      port map(A_DOUT(17) => nc151, A_DOUT(16) => nc23, 
        A_DOUT(15) => nc58, A_DOUT(14) => nc116, A_DOUT(13) => 
        nc74, A_DOUT(12) => nc133, A_DOUT(11) => nc167, 
        A_DOUT(10) => nc84, A_DOUT(9) => nc39, A_DOUT(8) => nc72, 
        A_DOUT(7) => nc82, A_DOUT(6) => nc145, A_DOUT(5) => nc160, 
        A_DOUT(4) => nc57, A_DOUT(3) => nc156, A_DOUT(2) => nc125, 
        A_DOUT(1) => RDATA_int(5), A_DOUT(0) => RDATA_int(4), 
        B_DOUT(17) => nc73, B_DOUT(16) => nc107, B_DOUT(15) => 
        nc66, B_DOUT(14) => nc83, B_DOUT(13) => nc9, B_DOUT(12)
         => nc171, B_DOUT(11) => nc54, B_DOUT(10) => nc135, 
        B_DOUT(9) => nc41, B_DOUT(8) => nc100, B_DOUT(7) => nc52, 
        B_DOUT(6) => nc29, B_DOUT(5) => nc118, B_DOUT(4) => nc60, 
        B_DOUT(3) => nc141, B_DOUT(2) => nc45, B_DOUT(1) => nc53, 
        B_DOUT(0) => nc121, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_283_i, A_BLK(1) => VCC_net_1, A_BLK(0) => VCC_net_1, 
        A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => VCC_net_1, 
        A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, A_DIN(15)
         => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13) => 
        GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => GND_net_1, 
        A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, A_DIN(8)
         => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6) => 
        GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => GND_net_1, 
        A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, A_DIN(1)
         => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13) => 
        fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(5), B_DIN(0) => RX_FIFO_DIN_pipe(4), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C1 : RAM1K18
      port map(A_DOUT(17) => nc158, A_DOUT(16) => nc162, 
        A_DOUT(15) => nc11, A_DOUT(14) => nc131, A_DOUT(13) => 
        nc96, A_DOUT(12) => nc79, A_DOUT(11) => nc146, A_DOUT(10)
         => nc89, A_DOUT(9) => nc119, A_DOUT(8) => nc48, 
        A_DOUT(7) => nc126, A_DOUT(6) => nc15, A_DOUT(5) => nc102, 
        A_DOUT(4) => nc3, A_DOUT(3) => nc47, A_DOUT(2) => nc90, 
        A_DOUT(1) => RDATA_int(3), A_DOUT(0) => RDATA_int(2), 
        B_DOUT(17) => nc159, B_DOUT(16) => nc136, B_DOUT(15) => 
        nc59, B_DOUT(14) => nc18, B_DOUT(13) => nc44, B_DOUT(12)
         => nc117, B_DOUT(11) => nc164, B_DOUT(10) => nc148, 
        B_DOUT(9) => nc42, B_DOUT(8) => nc17, B_DOUT(7) => nc2, 
        B_DOUT(6) => nc110, B_DOUT(5) => nc128, B_DOUT(4) => nc43, 
        B_DOUT(3) => nc157, B_DOUT(2) => nc36, B_DOUT(1) => nc61, 
        B_DOUT(0) => nc104, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_283_i, A_BLK(1) => VCC_net_1, A_BLK(0) => VCC_net_1, 
        A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => VCC_net_1, 
        A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, A_DIN(15)
         => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13) => 
        GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => GND_net_1, 
        A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, A_DIN(8)
         => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6) => 
        GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => GND_net_1, 
        A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, A_DIN(1)
         => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13) => 
        fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(3), B_DIN(0) => RX_FIFO_DIN_pipe(2), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C4 : RAM1K18
      port map(A_DOUT(17) => nc138, A_DOUT(16) => nc14, 
        A_DOUT(15) => nc150, A_DOUT(14) => nc149, A_DOUT(13) => 
        nc12, A_DOUT(12) => nc30, A_DOUT(11) => nc65, A_DOUT(10)
         => nc7, A_DOUT(9) => nc129, A_DOUT(8) => nc8, A_DOUT(7)
         => nc13, A_DOUT(6) => nc26, A_DOUT(5) => nc139, 
        A_DOUT(4) => nc163, A_DOUT(3) => nc112, A_DOUT(2) => nc68, 
        A_DOUT(1) => nc49, A_DOUT(0) => RDATA_int(8), B_DOUT(17)
         => nc170, B_DOUT(16) => nc91, B_DOUT(15) => nc5, 
        B_DOUT(14) => nc20, B_DOUT(13) => nc147, B_DOUT(12) => 
        nc67, B_DOUT(11) => nc152, B_DOUT(10) => nc127, B_DOUT(9)
         => nc103, B_DOUT(8) => nc76, B_DOUT(7) => nc140, 
        B_DOUT(6) => nc86, B_DOUT(5) => nc95, B_DOUT(4) => nc120, 
        B_DOUT(3) => nc165, B_DOUT(2) => nc137, B_DOUT(1) => nc64, 
        B_DOUT(0) => nc19, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_283_i, A_BLK(1) => VCC_net_1, A_BLK(0) => VCC_net_1, 
        A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => VCC_net_1, 
        A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, A_DIN(15)
         => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13) => 
        GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => GND_net_1, 
        A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, A_DIN(8)
         => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6) => 
        GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => GND_net_1, 
        A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, A_DIN(1)
         => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13) => 
        fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => GND_net_1, B_DIN(0) => RX_FIFO_DIN_pipe(8), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C3 : RAM1K18
      port map(A_DOUT(17) => nc70, A_DOUT(16) => nc62, A_DOUT(15)
         => nc80, A_DOUT(14) => nc130, A_DOUT(13) => nc98, 
        A_DOUT(12) => nc114, A_DOUT(11) => nc56, A_DOUT(10) => 
        nc105, A_DOUT(9) => nc63, A_DOUT(8) => nc97, A_DOUT(7)
         => nc161, A_DOUT(6) => nc31, A_DOUT(5) => nc154, 
        A_DOUT(4) => nc50, A_DOUT(3) => nc142, A_DOUT(2) => nc94, 
        A_DOUT(1) => RDATA_int(7), A_DOUT(0) => RDATA_int(6), 
        B_DOUT(17) => nc122, B_DOUT(16) => nc35, B_DOUT(15) => 
        nc4, B_DOUT(14) => nc92, B_DOUT(13) => nc101, B_DOUT(12)
         => nc166, B_DOUT(11) => nc132, B_DOUT(10) => nc21, 
        B_DOUT(9) => nc93, B_DOUT(8) => nc69, B_DOUT(7) => nc38, 
        B_DOUT(6) => nc113, B_DOUT(5) => nc106, B_DOUT(4) => nc25, 
        B_DOUT(3) => nc1, B_DOUT(2) => nc37, B_DOUT(1) => nc144, 
        B_DOUT(0) => nc153, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_283_i, A_BLK(1) => VCC_net_1, A_BLK(0) => VCC_net_1, 
        A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => VCC_net_1, 
        A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, A_DIN(15)
         => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13) => 
        GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => GND_net_1, 
        A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, A_DIN(8)
         => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6) => 
        GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => GND_net_1, 
        A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, A_DIN(1)
         => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13) => 
        fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(7), B_DIN(0) => RX_FIFO_DIN_pipe(6), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C0 : RAM1K18
      port map(A_DOUT(17) => nc46, A_DOUT(16) => nc71, A_DOUT(15)
         => nc124, A_DOUT(14) => nc81, A_DOUT(13) => nc168, 
        A_DOUT(12) => nc34, A_DOUT(11) => nc28, A_DOUT(10) => 
        nc115, A_DOUT(9) => nc134, A_DOUT(8) => nc32, A_DOUT(7)
         => nc40, A_DOUT(6) => nc99, A_DOUT(5) => nc75, A_DOUT(4)
         => nc85, A_DOUT(3) => nc27, A_DOUT(2) => nc108, 
        A_DOUT(1) => RDATA_int(1), A_DOUT(0) => RDATA_int(0), 
        B_DOUT(17) => nc16, B_DOUT(16) => nc155, B_DOUT(15) => 
        nc51, B_DOUT(14) => nc33, B_DOUT(13) => nc169, B_DOUT(12)
         => nc78, B_DOUT(11) => nc24, B_DOUT(10) => nc88, 
        B_DOUT(9) => nc111, B_DOUT(8) => nc55, B_DOUT(7) => nc10, 
        B_DOUT(6) => nc22, B_DOUT(5) => nc143, B_DOUT(4) => nc77, 
        B_DOUT(3) => nc6, B_DOUT(2) => nc109, B_DOUT(1) => nc87, 
        B_DOUT(0) => nc123, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_283_i, A_BLK(1) => VCC_net_1, A_BLK(0) => VCC_net_1, 
        A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => VCC_net_1, 
        A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, A_DIN(15)
         => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13) => 
        GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => GND_net_1, 
        A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, A_DIN(8)
         => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6) => 
        GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => GND_net_1, 
        A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, A_DIN(1)
         => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13) => 
        fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(1), B_DIN(0) => RX_FIFO_DIN_pipe(0), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper is

    port( fifo_MEMRADDR             : in    std_logic_vector(12 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0);
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          N_283_i                   : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          fifo_MEMWE                : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top
    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          fifo_MEMRADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          fifo_MEMWE                : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          N_283_i                   : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    L1_asyncnonpipe : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top
      port map(RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), RDATA_int(8)
         => RDATA_int(8), RDATA_int(7) => RDATA_int(7), 
        RDATA_int(6) => RDATA_int(6), RDATA_int(5) => 
        RDATA_int(5), RDATA_int(4) => RDATA_int(4), RDATA_int(3)
         => RDATA_int(3), RDATA_int(2) => RDATA_int(2), 
        RDATA_int(1) => RDATA_int(1), RDATA_int(0) => 
        RDATA_int(0), fifo_MEMWADDR(12) => fifo_MEMWADDR(12), 
        fifo_MEMWADDR(11) => fifo_MEMWADDR(11), fifo_MEMWADDR(10)
         => fifo_MEMWADDR(10), fifo_MEMWADDR(9) => 
        fifo_MEMWADDR(9), fifo_MEMWADDR(8) => fifo_MEMWADDR(8), 
        fifo_MEMWADDR(7) => fifo_MEMWADDR(7), fifo_MEMWADDR(6)
         => fifo_MEMWADDR(6), fifo_MEMWADDR(5) => 
        fifo_MEMWADDR(5), fifo_MEMWADDR(4) => fifo_MEMWADDR(4), 
        fifo_MEMWADDR(3) => fifo_MEMWADDR(3), fifo_MEMWADDR(2)
         => fifo_MEMWADDR(2), fifo_MEMWADDR(1) => 
        fifo_MEMWADDR(1), fifo_MEMWADDR(0) => fifo_MEMWADDR(0), 
        fifo_MEMRADDR(12) => fifo_MEMRADDR(12), fifo_MEMRADDR(11)
         => fifo_MEMRADDR(11), fifo_MEMRADDR(10) => 
        fifo_MEMRADDR(10), fifo_MEMRADDR(9) => fifo_MEMRADDR(9), 
        fifo_MEMRADDR(8) => fifo_MEMRADDR(8), fifo_MEMRADDR(7)
         => fifo_MEMRADDR(7), fifo_MEMRADDR(6) => 
        fifo_MEMRADDR(6), fifo_MEMRADDR(5) => fifo_MEMRADDR(5), 
        fifo_MEMRADDR(4) => fifo_MEMRADDR(4), fifo_MEMRADDR(3)
         => fifo_MEMRADDR(3), fifo_MEMRADDR(2) => 
        fifo_MEMRADDR(2), fifo_MEMRADDR(1) => fifo_MEMRADDR(1), 
        fifo_MEMRADDR(0) => fifo_MEMRADDR(0), fifo_MEMWE => 
        fifo_MEMWE, CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        N_283_i => N_283_i, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_0 is

    port( wptr_bin_sync  : inout std_logic_vector(13 downto 0) := (others => 'Z');
          wptr_gray_sync : in    std_logic_vector(12 downto 0);
          bin_N_6_i      : out   std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_0;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \bin_m5_5\, \bin_m5_4\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    bin_m5_4 : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(5), B => wptr_gray_sync(6), C
         => wptr_gray_sync(4), D => wptr_gray_sync(7), Y => 
        \bin_m5_4\);
    
    \bin_out_xhdl1_0_a2[10]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(12), B => wptr_bin_sync(13), C
         => wptr_gray_sync(10), D => wptr_gray_sync(11), Y => 
        wptr_bin_sync(10));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(8), B => wptr_gray_sync(9), C
         => wptr_bin_sync(10), Y => wptr_bin_sync(8));
    
    bin_m5_5 : CFG4
      generic map(INIT => x"9669")

      port map(A => wptr_gray_sync(10), B => wptr_gray_sync(11), 
        C => wptr_gray_sync(8), D => wptr_gray_sync(9), Y => 
        \bin_m5_5\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(3), B => wptr_gray_sync(2), Y
         => wptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[1]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(1), B => wptr_gray_sync(2), C
         => wptr_bin_sync(3), Y => wptr_bin_sync(1));
    
    \bin_out_xhdl1_i_o2_RNIKRPL2[12]\ : CFG3
      generic map(INIT => x"69")

      port map(A => \bin_m5_5\, B => \bin_m5_4\, C => 
        wptr_bin_sync(12), Y => bin_N_6_i);
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(1), B => wptr_gray_sync(0), C
         => wptr_bin_sync(3), D => wptr_gray_sync(2), Y => 
        wptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2[11]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(11), B => wptr_bin_sync(13), C
         => wptr_gray_sync(12), Y => wptr_bin_sync(11));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(9), B => wptr_bin_sync(10), C
         => wptr_gray_sync(7), D => wptr_gray_sync(8), Y => 
        wptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[5]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(5), B => wptr_gray_sync(6), C
         => wptr_bin_sync(7), Y => wptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(7), B => wptr_gray_sync(6), Y
         => wptr_bin_sync(6));
    
    \bin_out_xhdl1_i_o2[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(13), B => wptr_gray_sync(12), Y
         => wptr_bin_sync(12));
    
    \bin_out_xhdl1_0_a2[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(10), B => wptr_gray_sync(9), Y
         => wptr_bin_sync(9));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"9669")

      port map(A => wptr_bin_sync(12), B => \bin_m5_5\, C => 
        wptr_gray_sync(3), D => \bin_m5_4\, Y => wptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1 is

    port( wptr_gray                 : in    std_logic_vector(13 downto 0);
          wptr_gray_sync            : out   std_logic_vector(12 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \sync_int[11]_net_1\, GND_net_1, 
        \sync_int[12]_net_1\, \sync_int[13]_net_1\, 
        \sync_int[10]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\, \sync_int[4]_net_1\, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => wptr_gray(9), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => wptr_gray(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => wptr_gray(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => wptr_gray(11), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => wptr_gray(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(11));
    
    \sync_int[13]\ : SLE
      port map(D => wptr_gray(13), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[13]_net_1\);
    
    \sync_int[3]\ : SLE
      port map(D => wptr_gray(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[3]_net_1\);
    
    \sync_int[12]\ : SLE
      port map(D => wptr_gray(12), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[12]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => wptr_gray(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => wptr_gray(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => wptr_gray(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[12]\ : SLE
      port map(D => \sync_int[12]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(12));
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => wptr_gray(8), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => wptr_gray(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => wptr_gray(10), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[10]_net_1\);
    
    \sync_out_xhdl1[13]\ : SLE
      port map(D => \sync_int[13]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_bin_sync_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0 is

    port( rptr_gray           : in    std_logic_vector(13 downto 0);
          rptr_gray_sync      : out   std_logic_vector(12 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          irx_fifo_rst_i      : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \sync_int[13]_net_1\, GND_net_1, 
        \sync_int[12]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\, \sync_int[4]_net_1\, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\, \sync_int[10]_net_1\, 
        \sync_int[11]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => rptr_gray(9), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => rptr_gray(4), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => rptr_gray(1), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => rptr_gray(11), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => rptr_gray(6), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(11));
    
    \sync_int[13]\ : SLE
      port map(D => rptr_gray(13), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[13]_net_1\);
    
    \sync_int[3]\ : SLE
      port map(D => rptr_gray(3), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[3]_net_1\);
    
    \sync_int[12]\ : SLE
      port map(D => rptr_gray(12), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[12]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => rptr_gray(0), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => rptr_gray(5), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => rptr_gray(2), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[12]\ : SLE
      port map(D => \sync_int[12]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(12));
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => rptr_gray(8), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => rptr_gray(7), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => rptr_gray(10), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[10]_net_1\);
    
    \sync_out_xhdl1[13]\ : SLE
      port map(D => \sync_int[13]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_bin_sync_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv is

    port( rptr_bin_sync  : inout std_logic_vector(13 downto 0) := (others => 'Z');
          rptr_gray_sync : in    std_logic_vector(12 downto 0);
          bin_N_6_i      : out   std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \bin_m5_5\, \bin_m5_4\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    bin_m5_4 : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(5), B => rptr_gray_sync(6), C
         => rptr_gray_sync(4), D => rptr_gray_sync(7), Y => 
        \bin_m5_4\);
    
    \bin_out_xhdl1_i_o2_RNI99AG2[12]\ : CFG3
      generic map(INIT => x"69")

      port map(A => \bin_m5_5\, B => \bin_m5_4\, C => 
        rptr_bin_sync(12), Y => bin_N_6_i);
    
    \bin_out_xhdl1_0_a2[10]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(12), B => rptr_bin_sync(13), C
         => rptr_gray_sync(10), D => rptr_gray_sync(11), Y => 
        rptr_bin_sync(10));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(8), B => rptr_gray_sync(9), C
         => rptr_bin_sync(10), Y => rptr_bin_sync(8));
    
    bin_m5_5 : CFG4
      generic map(INIT => x"9669")

      port map(A => rptr_gray_sync(10), B => rptr_gray_sync(11), 
        C => rptr_gray_sync(8), D => rptr_gray_sync(9), Y => 
        \bin_m5_5\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(3), B => rptr_gray_sync(2), Y
         => rptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[1]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(1), B => rptr_gray_sync(2), C
         => rptr_bin_sync(3), Y => rptr_bin_sync(1));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(1), B => rptr_gray_sync(0), C
         => rptr_bin_sync(3), D => rptr_gray_sync(2), Y => 
        rptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2[11]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(11), B => rptr_bin_sync(13), C
         => rptr_gray_sync(12), Y => rptr_bin_sync(11));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(8), B => rptr_gray_sync(7), C
         => rptr_bin_sync(10), D => rptr_gray_sync(9), Y => 
        rptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[5]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(5), B => rptr_gray_sync(6), C
         => rptr_bin_sync(7), Y => rptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(7), B => rptr_gray_sync(6), Y
         => rptr_bin_sync(6));
    
    \bin_out_xhdl1_i_o2[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(13), B => rptr_gray_sync(12), Y
         => rptr_bin_sync(12));
    
    \bin_out_xhdl1_0_a2[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(10), B => rptr_gray_sync(9), Y
         => rptr_bin_sync(9));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"9669")

      port map(A => rptr_bin_sync(12), B => \bin_m5_5\, C => 
        rptr_gray_sync(3), D => \bin_m5_4\, Y => rptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async is

    port( rdiff_bus                 : out   std_logic_vector(13 downto 1);
          fifo_MEMRADDR             : out   std_logic_vector(12 downto 0);
          fifo_MEMWADDR             : out   std_logic_vector(12 downto 0);
          tx_col_detect_en          : in    std_logic;
          RX_InProcess_d1           : in    std_logic;
          sampler_clk1x_en          : in    std_logic;
          iRX_FIFO_wr_en            : in    std_logic;
          rdiff_bus_cry_0_Y_0       : out   std_logic;
          un2_re_p                  : in    std_logic;
          RX_FIFO_Full              : out   std_logic;
          empty_r_3                 : in    std_logic;
          RX_FIFO_Empty             : out   std_logic;
          N_283_i                   : in    std_logic;
          fifo_MEMWE                : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          irx_fifo_rst_i            : in    std_logic;
          RX_FIFO_OVERFLOW_i        : out   std_logic;
          RX_FIFO_OVERFLOW          : out   std_logic;
          RX_FIFO_UNDERRUN_i        : out   std_logic;
          RX_FIFO_UNDERRUN          : out   std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_0
    port( wptr_bin_sync  : inout   std_logic_vector(13 downto 0);
          wptr_gray_sync : in    std_logic_vector(12 downto 0) := (others => 'U');
          bin_N_6_i      : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1
    port( wptr_gray                 : in    std_logic_vector(13 downto 0) := (others => 'U');
          wptr_gray_sync            : out   std_logic_vector(12 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0
    port( rptr_gray           : in    std_logic_vector(13 downto 0) := (others => 'U');
          rptr_gray_sync      : out   std_logic_vector(12 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          irx_fifo_rst_i      : in    std_logic := 'U'
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv
    port( rptr_bin_sync  : inout   std_logic_vector(13 downto 0);
          rptr_gray_sync : in    std_logic_vector(12 downto 0) := (others => 'U');
          bin_N_6_i      : out   std_logic
        );
  end component;

    signal \rptr[0]_net_1\, \rptr_s[0]\, \fifo_MEMRADDR[0]\, 
        \fifo_MEMRADDR_i[0]\, \fifo_MEMWADDR[0]\, 
        \fifo_MEMWADDR_i[0]\, \RX_FIFO_UNDERRUN\, 
        \RX_FIFO_OVERFLOW\, \wptr_gray[1]_net_1\, VCC_net_1, 
        \wptr_gray_1[1]_net_1\, GND_net_1, \wptr_gray[2]_net_1\, 
        \wptr_gray_1[2]_net_1\, \wptr_gray[3]_net_1\, 
        \wptr_gray_1[3]_net_1\, \wptr_gray[4]_net_1\, 
        \wptr_gray_1[4]_net_1\, \wptr_gray[5]_net_1\, 
        \wptr_gray_1[5]_net_1\, \wptr_gray[6]_net_1\, 
        \wptr_gray_1[6]_net_1\, \wptr_gray[7]_net_1\, 
        \wptr_gray_1[7]_net_1\, \wptr_gray[8]_net_1\, 
        \wptr_gray_1[8]_net_1\, \wptr_gray[9]_net_1\, 
        \wptr_gray_1[9]_net_1\, \wptr_gray[10]_net_1\, 
        \wptr_gray_1[10]_net_1\, \wptr_gray[11]_net_1\, 
        \wptr_gray_1[11]_net_1\, \wptr_gray[12]_net_1\, 
        \wptr_gray_1[12]_net_1\, \wptr_gray[13]_net_1\, 
        \wptr[13]_net_1\, \rptr_bin_sync2[0]_net_1\, 
        \rptr_bin_sync[0]\, \rptr_bin_sync2[1]_net_1\, 
        \rptr_bin_sync[1]\, \rptr_bin_sync2[2]_net_1\, 
        \rptr_bin_sync[2]\, \rptr_bin_sync2[3]_net_1\, 
        \rptr_bin_sync[3]\, \rptr_bin_sync2[4]_net_1\, bin_N_6_i, 
        \rptr_bin_sync2[5]_net_1\, \rptr_bin_sync[5]\, 
        \rptr_bin_sync2[6]_net_1\, \rptr_bin_sync[6]\, 
        \rptr_bin_sync2[7]_net_1\, \rptr_bin_sync[7]\, 
        \rptr_bin_sync2[8]_net_1\, \rptr_bin_sync[8]\, 
        \rptr_bin_sync2[9]_net_1\, \rptr_bin_sync[9]\, 
        \rptr_bin_sync2[10]_net_1\, \rptr_bin_sync[10]\, 
        \rptr_bin_sync2[11]_net_1\, \rptr_bin_sync[11]\, 
        \rptr_bin_sync2[12]_net_1\, \rptr_bin_sync[12]\, 
        \rptr_bin_sync2[13]_net_1\, \rptr_bin_sync[13]\, 
        \wptr_gray[0]_net_1\, \wptr_gray_1[0]_net_1\, \rdiff_bus\, 
        \wptr_bin_sync[0]\, \wptr_bin_sync2[1]_net_1\, 
        \wptr_bin_sync[1]\, \wptr_bin_sync2[2]_net_1\, 
        \wptr_bin_sync[2]\, \wptr_bin_sync2[3]_net_1\, 
        \wptr_bin_sync[3]\, \wptr_bin_sync2[4]_net_1\, 
        bin_N_6_i_0, \wptr_bin_sync2[5]_net_1\, 
        \wptr_bin_sync[5]\, \wptr_bin_sync2[6]_net_1\, 
        \wptr_bin_sync[6]\, \wptr_bin_sync2[7]_net_1\, 
        \wptr_bin_sync[7]\, \wptr_bin_sync2[8]_net_1\, 
        \wptr_bin_sync[8]\, \wptr_bin_sync2[9]_net_1\, 
        \wptr_bin_sync[9]\, \wptr_bin_sync2[10]_net_1\, 
        \wptr_bin_sync[10]\, \wptr_bin_sync2[11]_net_1\, 
        \wptr_bin_sync[11]\, \wptr_bin_sync2[12]_net_1\, 
        \wptr_bin_sync[12]\, \wptr_bin_sync2[13]_net_1\, 
        \wptr_bin_sync[13]\, \rptr_gray[9]_net_1\, 
        \rptr_gray_1[9]_net_1\, \rptr_gray[10]_net_1\, 
        \rptr_gray_1[10]_net_1\, \rptr_gray[11]_net_1\, 
        \rptr_gray_1[11]_net_1\, \rptr_gray[12]_net_1\, 
        \rptr_gray_1[12]_net_1\, \rptr_gray[13]_net_1\, 
        \rptr[13]_net_1\, \fifo_MEMWADDR[7]\, 
        \memwaddr_r_2[7]_net_1\, \fifo_MEMWE\, \fifo_MEMWADDR[8]\, 
        \memwaddr_r_2[8]_net_1\, \fifo_MEMWADDR[9]\, 
        \memwaddr_r_2[9]_net_1\, \fifo_MEMWADDR[10]\, 
        \memwaddr_r_2[10]_net_1\, \fifo_MEMWADDR[11]\, 
        \memwaddr_r_2[11]_net_1\, \fifo_MEMWADDR[12]\, 
        \memwaddr_r_2[12]_net_1\, \rptr_gray[0]_net_1\, 
        \rptr_gray_1[0]_net_1\, \rptr_gray[1]_net_1\, 
        \rptr_gray_1[1]_net_1\, \rptr_gray[2]_net_1\, 
        \rptr_gray_1[2]_net_1\, \rptr_gray[3]_net_1\, 
        \rptr_gray_1[3]_net_1\, \rptr_gray[4]_net_1\, 
        \rptr_gray_1[4]_net_1\, \rptr_gray[5]_net_1\, 
        \rptr_gray_1[5]_net_1\, \rptr_gray[6]_net_1\, 
        \rptr_gray_1[6]_net_1\, \rptr_gray[7]_net_1\, 
        \rptr_gray_1[7]_net_1\, \rptr_gray[8]_net_1\, 
        \rptr_gray_1[8]_net_1\, \fifo_MEMRADDR[5]\, 
        \memraddr_r_2[5]_net_1\, \fifo_MEMRADDR[6]\, 
        un1_memraddr_r_cry_6_S, \fifo_MEMRADDR[7]\, 
        \memraddr_r_2[7]_net_1\, \fifo_MEMRADDR[8]\, 
        \memraddr_r_2[8]_net_1\, \fifo_MEMRADDR[9]\, 
        \memraddr_r_2[9]_net_1\, \fifo_MEMRADDR[10]\, 
        \memraddr_r_2[10]_net_1\, \fifo_MEMRADDR[11]\, 
        \memraddr_r_2[11]_net_1\, \fifo_MEMRADDR[12]\, 
        \memraddr_r_2[12]_net_1\, \fifo_MEMWADDR[1]\, 
        un1_memwaddr_r_cry_1_S, \fifo_MEMWADDR[2]\, 
        un1_memwaddr_r_cry_2_S, \fifo_MEMWADDR[3]\, 
        un1_memwaddr_r_cry_3_S, \fifo_MEMWADDR[4]\, 
        un1_memwaddr_r_cry_4_S, \fifo_MEMWADDR[5]\, 
        \memwaddr_r_2[5]_net_1\, \fifo_MEMWADDR[6]\, 
        un1_memwaddr_r_cry_6_S, \fifo_MEMRADDR[1]\, 
        un1_memraddr_r_cry_1_S, \fifo_MEMRADDR[2]\, 
        un1_memraddr_r_cry_2_S, \fifo_MEMRADDR[3]\, 
        un1_memraddr_r_cry_3_S, \fifo_MEMRADDR[4]\, 
        un1_memraddr_r_cry_4_S, \RX_FIFO_Full\, fulli, un1_we_p, 
        \rptr[1]_net_1\, \rptr_s[1]\, \rptr[2]_net_1\, 
        \rptr_s[2]\, \rptr[3]_net_1\, \rptr_s[3]\, 
        \rptr[4]_net_1\, \rptr_s[4]\, \rptr[5]_net_1\, 
        \rptr_s[5]\, \rptr[6]_net_1\, \rptr_s[6]\, 
        \rptr[7]_net_1\, \rptr_s[7]\, \rptr[8]_net_1\, 
        \rptr_s[8]\, \rptr[9]_net_1\, \rptr_s[9]\, 
        \rptr[10]_net_1\, \rptr_s[10]\, \rptr[11]_net_1\, 
        \rptr_s[11]\, \rptr[12]_net_1\, \rptr_s[12]\, 
        \rptr_s[13]_net_1\, \wptr[0]_net_1\, \wptr_s[0]\, N_586, 
        \wptr[1]_net_1\, \wptr_s[1]\, \wptr[2]_net_1\, 
        \wptr_s[2]\, \wptr[3]_net_1\, \wptr_s[3]\, 
        \wptr[4]_net_1\, \wptr_s[4]\, \wptr[5]_net_1\, 
        \wptr_s[5]\, \wptr[6]_net_1\, \wptr_s[6]\, 
        \wptr[7]_net_1\, \wptr_s[7]\, \wptr[8]_net_1\, 
        \wptr_s[8]\, \wptr[9]_net_1\, \wptr_s[9]\, 
        \wptr[10]_net_1\, \wptr_s[10]\, \wptr[11]_net_1\, 
        \wptr_s[11]\, \wptr[12]_net_1\, \wptr_s[12]\, 
        \wptr_s[13]_net_1\, wptr_cry_cy, \wptr_cry[0]_net_1\, 
        \wptr_cry[1]_net_1\, \wptr_cry[2]_net_1\, 
        \wptr_cry[3]_net_1\, \wptr_cry[4]_net_1\, 
        \wptr_cry[5]_net_1\, \wptr_cry[6]_net_1\, 
        \wptr_cry[7]_net_1\, \wptr_cry[8]_net_1\, 
        \wptr_cry[9]_net_1\, \wptr_cry[10]_net_1\, 
        \wptr_cry[11]_net_1\, \wptr_cry[12]_net_1\, 
        \wdiff_bus_cry_0\, wdiff_bus_cry_0_Y_0, \wdiff_bus_cry_1\, 
        \wdiff_bus[1]\, \wdiff_bus_cry_2\, \wdiff_bus[2]\, 
        \wdiff_bus_cry_3\, \wdiff_bus[3]\, \wdiff_bus_cry_4\, 
        \wdiff_bus[4]\, \wdiff_bus_cry_5\, \wdiff_bus[5]\, 
        \wdiff_bus_cry_6\, \wdiff_bus[6]\, \wdiff_bus_cry_7\, 
        \wdiff_bus[7]\, \wdiff_bus_cry_8\, \wdiff_bus[8]\, 
        \wdiff_bus_cry_9\, \wdiff_bus[9]\, \wdiff_bus_cry_10\, 
        \wdiff_bus[10]\, \wdiff_bus_cry_11\, \wdiff_bus[11]\, 
        \wdiff_bus[13]\, \wdiff_bus_cry_12\, \wdiff_bus[12]\, 
        \rdiff_bus_cry_0\, \rdiff_bus_cry_1\, \rdiff_bus_cry_2\, 
        \rdiff_bus_cry_3\, \rdiff_bus_cry_4\, \rdiff_bus_cry_5\, 
        \rdiff_bus_cry_6\, \rdiff_bus_cry_7\, \rdiff_bus_cry_8\, 
        \rdiff_bus_cry_9\, \rdiff_bus_cry_10\, \rdiff_bus_cry_11\, 
        \rdiff_bus_cry_12\, rptr_s_266_FCO, \rptr_cry[1]_net_1\, 
        \rptr_cry[2]_net_1\, \rptr_cry[3]_net_1\, 
        \rptr_cry[4]_net_1\, \rptr_cry[5]_net_1\, 
        \rptr_cry[6]_net_1\, \rptr_cry[7]_net_1\, 
        \rptr_cry[8]_net_1\, \rptr_cry[9]_net_1\, 
        \rptr_cry[10]_net_1\, \rptr_cry[11]_net_1\, 
        \rptr_cry[12]_net_1\, un1_memraddr_r_s_1_275_FCO, 
        \un1_memraddr_r_cry_1\, \un1_memraddr_r_cry_2\, 
        \un1_memraddr_r_cry_3\, \un1_memraddr_r_cry_4\, 
        \un1_memraddr_r_cry_5\, un1_memraddr_r_cry_5_S, 
        \un1_memraddr_r_cry_6\, \un1_memraddr_r_cry_7\, 
        un1_memraddr_r_cry_7_S, \un1_memraddr_r_cry_8\, 
        un1_memraddr_r_cry_8_S, \un1_memraddr_r_cry_9\, 
        un1_memraddr_r_cry_9_S, \un1_memraddr_r_cry_10\, 
        un1_memraddr_r_cry_10_S, un1_memraddr_r_s_12_S, 
        \un1_memraddr_r_cry_11\, un1_memraddr_r_cry_11_S, 
        un1_memwaddr_r_s_1_276_FCO, \un1_memwaddr_r_cry_1\, 
        \un1_memwaddr_r_cry_2\, \un1_memwaddr_r_cry_3\, 
        \un1_memwaddr_r_cry_4\, \un1_memwaddr_r_cry_5\, 
        un1_memwaddr_r_cry_5_S, \un1_memwaddr_r_cry_6\, 
        \un1_memwaddr_r_cry_7\, un1_memwaddr_r_cry_7_S, 
        \un1_memwaddr_r_cry_8\, un1_memwaddr_r_cry_8_S, 
        \un1_memwaddr_r_cry_9\, un1_memwaddr_r_cry_9_S, 
        \un1_memwaddr_r_cry_10\, un1_memwaddr_r_cry_10_S, 
        un1_memwaddr_r_s_12_S, \un1_memwaddr_r_cry_11\, 
        un1_memwaddr_r_cry_11_S, \fulli_0_1\, \fulli_0_a2_3\, 
        N_567, un4_re_i_0, un4_we_i_0, un4_re_i_8, un4_re_i_7, 
        un4_we_i_8, un4_we_i_7, \fulli_0_a2_0_2\, un4_re_i_9, 
        un4_we_i_9, \wptr_gray_sync[0]\, \wptr_gray_sync[1]\, 
        \wptr_gray_sync[2]\, \wptr_gray_sync[3]\, 
        \wptr_gray_sync[4]\, \wptr_gray_sync[5]\, 
        \wptr_gray_sync[6]\, \wptr_gray_sync[7]\, 
        \wptr_gray_sync[8]\, \wptr_gray_sync[9]\, 
        \wptr_gray_sync[10]\, \wptr_gray_sync[11]\, 
        \wptr_gray_sync[12]\, \rptr_gray_sync[0]\, 
        \rptr_gray_sync[1]\, \rptr_gray_sync[2]\, 
        \rptr_gray_sync[3]\, \rptr_gray_sync[4]\, 
        \rptr_gray_sync[5]\, \rptr_gray_sync[6]\, 
        \rptr_gray_sync[7]\, \rptr_gray_sync[8]\, 
        \rptr_gray_sync[9]\, \rptr_gray_sync[10]\, 
        \rptr_gray_sync[11]\, \rptr_gray_sync[12]\ : std_logic;
    signal nc2, nc1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_0
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_0(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv(DEF_ARCH);
begin 

    fifo_MEMRADDR(12) <= \fifo_MEMRADDR[12]\;
    fifo_MEMRADDR(11) <= \fifo_MEMRADDR[11]\;
    fifo_MEMRADDR(10) <= \fifo_MEMRADDR[10]\;
    fifo_MEMRADDR(9) <= \fifo_MEMRADDR[9]\;
    fifo_MEMRADDR(8) <= \fifo_MEMRADDR[8]\;
    fifo_MEMRADDR(7) <= \fifo_MEMRADDR[7]\;
    fifo_MEMRADDR(6) <= \fifo_MEMRADDR[6]\;
    fifo_MEMRADDR(5) <= \fifo_MEMRADDR[5]\;
    fifo_MEMRADDR(4) <= \fifo_MEMRADDR[4]\;
    fifo_MEMRADDR(3) <= \fifo_MEMRADDR[3]\;
    fifo_MEMRADDR(2) <= \fifo_MEMRADDR[2]\;
    fifo_MEMRADDR(1) <= \fifo_MEMRADDR[1]\;
    fifo_MEMRADDR(0) <= \fifo_MEMRADDR[0]\;
    fifo_MEMWADDR(12) <= \fifo_MEMWADDR[12]\;
    fifo_MEMWADDR(11) <= \fifo_MEMWADDR[11]\;
    fifo_MEMWADDR(10) <= \fifo_MEMWADDR[10]\;
    fifo_MEMWADDR(9) <= \fifo_MEMWADDR[9]\;
    fifo_MEMWADDR(8) <= \fifo_MEMWADDR[8]\;
    fifo_MEMWADDR(7) <= \fifo_MEMWADDR[7]\;
    fifo_MEMWADDR(6) <= \fifo_MEMWADDR[6]\;
    fifo_MEMWADDR(5) <= \fifo_MEMWADDR[5]\;
    fifo_MEMWADDR(4) <= \fifo_MEMWADDR[4]\;
    fifo_MEMWADDR(3) <= \fifo_MEMWADDR[3]\;
    fifo_MEMWADDR(2) <= \fifo_MEMWADDR[2]\;
    fifo_MEMWADDR(1) <= \fifo_MEMWADDR[1]\;
    fifo_MEMWADDR(0) <= \fifo_MEMWADDR[0]\;
    RX_FIFO_Full <= \RX_FIFO_Full\;
    fifo_MEMWE <= \fifo_MEMWE\;
    RX_FIFO_OVERFLOW <= \RX_FIFO_OVERFLOW\;
    RX_FIFO_UNDERRUN <= \RX_FIFO_UNDERRUN\;

    \rptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[4]_net_1\, S
         => \rptr_s[5]\, Y => OPEN, FCO => \rptr_cry[5]_net_1\);
    
    \memwaddr_r_2[9]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_9_S, D => un4_we_i_9, Y => 
        \memwaddr_r_2[9]_net_1\);
    
    wdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[8]_net_1\, B => 
        \rptr_bin_sync2[8]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_7\, S => \wdiff_bus[8]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_8\);
    
    \wptr_bin_sync2[12]\ : SLE
      port map(D => \wptr_bin_sync[12]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[12]_net_1\);
    
    wdiff_bus_cry_11 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[11]_net_1\, B => 
        \rptr_bin_sync2[11]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_10\, S => 
        \wdiff_bus[11]\, Y => OPEN, FCO => \wdiff_bus_cry_11\);
    
    un1_memwaddr_r_s_1_276 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => un1_memwaddr_r_s_1_276_FCO);
    
    \wptr_gray[4]\ : SLE
      port map(D => \wptr_gray_1[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[4]_net_1\);
    
    \rptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[3]_net_1\, B => \rptr[4]_net_1\, Y => 
        \rptr_gray_1[3]_net_1\);
    
    \rptr_bin_sync2[6]\ : SLE
      port map(D => \rptr_bin_sync[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[6]_net_1\);
    
    \rptr[1]\ : SLE
      port map(D => \rptr_s[1]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => N_283_i, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[1]_net_1\);
    
    \wptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[9]_net_1\, B => \wptr[10]_net_1\, Y => 
        \wptr_gray_1[9]_net_1\);
    
    \rptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[5]_net_1\, B => \rptr[6]_net_1\, Y => 
        \rptr_gray_1[5]_net_1\);
    
    \rptr_gray[9]\ : SLE
      port map(D => \rptr_gray_1[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[9]_net_1\);
    
    un1_memwaddr_r_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_6\, 
        S => un1_memwaddr_r_cry_7_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_7\);
    
    \rptr_gray[8]\ : SLE
      port map(D => \rptr_gray_1[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[8]_net_1\);
    
    un1_memraddr_r_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[11]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_10\, 
        S => un1_memraddr_r_cry_11_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_11\);
    
    \rptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[2]_net_1\, B => \rptr[3]_net_1\, Y => 
        \rptr_gray_1[2]_net_1\);
    
    \rptr_bin_sync2[7]\ : SLE
      port map(D => \rptr_bin_sync[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[7]_net_1\);
    
    \memwaddr_r[1]\ : SLE
      port map(D => un1_memwaddr_r_cry_1_S, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[1]\);
    
    rptr_s_266 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => rptr_s_266_FCO);
    
    \wptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[7]_net_1\, B => \wptr[8]_net_1\, Y => 
        \wptr_gray_1[7]_net_1\);
    
    \rptr_gray[13]\ : SLE
      port map(D => \rptr[13]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[13]_net_1\);
    
    \memraddr_r[0]\ : SLE
      port map(D => \fifo_MEMRADDR_i[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_283_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[0]\);
    
    \memraddr_r_2[9]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_9_S, D => un4_re_i_9, Y => 
        \memraddr_r_2[9]_net_1\);
    
    \wptr[0]\ : SLE
      port map(D => \wptr_s[0]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => N_586, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr[0]_net_1\);
    
    \rptr_bin_sync2[8]\ : SLE
      port map(D => \rptr_bin_sync[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[8]_net_1\);
    
    \rptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[1]_net_1\, B => \rptr[2]_net_1\, Y => 
        \rptr_gray_1[1]_net_1\);
    
    \rptr_gray[10]\ : SLE
      port map(D => \rptr_gray_1[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[10]_net_1\);
    
    \wptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[1]_net_1\, B => \wptr[0]_net_1\, Y => 
        \wptr_gray_1[0]_net_1\);
    
    wdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[9]_net_1\, B => 
        \rptr_bin_sync2[9]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_8\, S => \wdiff_bus[9]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_9\);
    
    \rptr[5]\ : SLE
      port map(D => \rptr_s[5]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => N_283_i, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[5]_net_1\);
    
    \rptr_gray[3]\ : SLE
      port map(D => \rptr_gray_1[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[3]_net_1\);
    
    \rptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[5]_net_1\, S
         => \rptr_s[6]\, Y => OPEN, FCO => \rptr_cry[6]_net_1\);
    
    \wptr_gray[3]\ : SLE
      port map(D => \wptr_gray_1[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[3]_net_1\);
    
    \rptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[10]_net_1\, B => \rptr[11]_net_1\, Y
         => \rptr_gray_1[10]_net_1\);
    
    un1_memraddr_r_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_9\, 
        S => un1_memraddr_r_cry_10_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_10\);
    
    \rptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[7]_net_1\, S
         => \rptr_s[8]\, Y => OPEN, FCO => \rptr_cry[8]_net_1\);
    
    \rptr[7]\ : SLE
      port map(D => \rptr_s[7]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => N_283_i, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[7]_net_1\);
    
    rdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[4]_net_1\, B => 
        \rptr[4]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_3\, S => rdiff_bus(4), Y => OPEN, FCO => 
        \rdiff_bus_cry_4\);
    
    \rptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[9]_net_1\, S
         => \rptr_s[10]\, Y => OPEN, FCO => \rptr_cry[10]_net_1\);
    
    \rptr_bin_sync2[12]\ : SLE
      port map(D => \rptr_bin_sync[12]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[12]_net_1\);
    
    \rptr_bin_sync2[0]\ : SLE
      port map(D => \rptr_bin_sync[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[0]_net_1\);
    
    \wptr[11]\ : SLE
      port map(D => \wptr_s[11]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => N_586, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr[11]_net_1\);
    
    rdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[1]_net_1\, B => 
        \rptr[1]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_0\, S => rdiff_bus(1), Y => OPEN, FCO => 
        \rdiff_bus_cry_1\);
    
    \memraddr_r[1]\ : SLE
      port map(D => un1_memraddr_r_cry_1_S, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_283_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[1]\);
    
    \L1.un1_we_p_0_a2_0\ : CFG4
      generic map(INIT => x"0080")

      port map(A => iRX_FIFO_wr_en, B => sampler_clk1x_en, C => 
        RX_InProcess_d1, D => tx_col_detect_en, Y => N_586);
    
    \rptr_bin_sync2[2]\ : SLE
      port map(D => \rptr_bin_sync[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[2]_net_1\);
    
    \memraddr_r_2[7]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_7_S, D => un4_re_i_9, Y => 
        \memraddr_r_2[7]_net_1\);
    
    un1_memwaddr_r_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_5\, 
        S => un1_memwaddr_r_cry_6_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_6\);
    
    rdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[6]_net_1\, B => 
        \rptr[6]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_5\, S => rdiff_bus(6), Y => OPEN, FCO => 
        \rdiff_bus_cry_6\);
    
    \memwaddr_r_2[10]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_10_S, D => un4_we_i_9, Y => 
        \memwaddr_r_2[10]_net_1\);
    
    \memraddr_r_2[5]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_5_S, D => un4_re_i_9, Y => 
        \memraddr_r_2[5]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    un1_memwaddr_r_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_8\, 
        S => un1_memwaddr_r_cry_9_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_9\);
    
    \rptr_gray[1]\ : SLE
      port map(D => \rptr_gray_1[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[1]_net_1\);
    
    \memwaddr_r[7]\ : SLE
      port map(D => \memwaddr_r_2[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[7]\);
    
    \wptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[3]_net_1\, S
         => \wptr_s[4]\, Y => OPEN, FCO => \wptr_cry[4]_net_1\);
    
    \wptr_gray_1[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[13]_net_1\, B => \wptr[12]_net_1\, Y
         => \wptr_gray_1[12]_net_1\);
    
    \wptr[12]\ : SLE
      port map(D => \wptr_s[12]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => N_586, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr[12]_net_1\);
    
    \wptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[9]_net_1\, S
         => \wptr_s[10]\, Y => OPEN, FCO => \wptr_cry[10]_net_1\);
    
    wdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[5]_net_1\, B => 
        \rptr_bin_sync2[5]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_4\, S => \wdiff_bus[5]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_5\);
    
    \rptr_gray[12]\ : SLE
      port map(D => \rptr_gray_1[12]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[12]_net_1\);
    
    \memwaddr_r[4]\ : SLE
      port map(D => un1_memwaddr_r_cry_4_S, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[4]\);
    
    \wptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[1]_net_1\, S
         => \wptr_s[2]\, Y => OPEN, FCO => \wptr_cry[2]_net_1\);
    
    \memraddr_r_2[10]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_10_S, D => un4_re_i_9, Y => 
        \memraddr_r_2[10]_net_1\);
    
    rdiff_bus_cry_11 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[11]_net_1\, B => 
        \rptr[11]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_10\, S => rdiff_bus(11), Y => OPEN, FCO
         => \rdiff_bus_cry_11\);
    
    fulli_0_a2_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => N_586, B => \fulli_0_a2_0_2\, C => 
        \wdiff_bus[3]\, D => \wdiff_bus[2]\, Y => N_567);
    
    wdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[0]_net_1\, B => 
        \rptr_bin_sync2[0]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => VCC_net_1, S => OPEN, Y => wdiff_bus_cry_0_Y_0, 
        FCO => \wdiff_bus_cry_0\);
    
    \wptr[1]\ : SLE
      port map(D => \wptr_s[1]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => N_586, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr[1]_net_1\);
    
    \rptr_bin_sync2[4]\ : SLE
      port map(D => bin_N_6_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[4]_net_1\);
    
    \wptr_bin_sync2[6]\ : SLE
      port map(D => \wptr_bin_sync[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[6]_net_1\);
    
    underflow_r_RNI7E0F : CFG1
      generic map(INIT => "01")

      port map(A => \RX_FIFO_UNDERRUN\, Y => RX_FIFO_UNDERRUN_i);
    
    \rptr[3]\ : SLE
      port map(D => \rptr_s[3]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => N_283_i, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[3]_net_1\);
    
    \wptr_gray[13]\ : SLE
      port map(D => \wptr[13]_net_1\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr_gray[13]_net_1\);
    
    \wptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[2]_net_1\, S
         => \wptr_s[3]\, Y => OPEN, FCO => \wptr_cry[3]_net_1\);
    
    \rptr[6]\ : SLE
      port map(D => \rptr_s[6]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => N_283_i, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[6]_net_1\);
    
    rdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[8]_net_1\, B => 
        \rptr[8]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_7\, S => rdiff_bus(8), Y => OPEN, FCO => 
        \rdiff_bus_cry_8\);
    
    \wptr_gray[10]\ : SLE
      port map(D => \wptr_gray_1[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[10]_net_1\);
    
    rdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[7]_net_1\, B => 
        \rptr[7]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_6\, S => rdiff_bus(7), Y => OPEN, FCO => 
        \rdiff_bus_cry_7\);
    
    \wptr_bin_sync2[7]\ : SLE
      port map(D => \wptr_bin_sync[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[7]_net_1\);
    
    \rptr_gray_1[11]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[11]_net_1\, B => \rptr[12]_net_1\, Y
         => \rptr_gray_1[11]_net_1\);
    
    \rptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[8]_net_1\, S
         => \rptr_s[9]\, Y => OPEN, FCO => \rptr_cry[9]_net_1\);
    
    un1_memwaddr_r_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        un1_memwaddr_r_s_1_276_FCO, S => un1_memwaddr_r_cry_1_S, 
        Y => OPEN, FCO => \un1_memwaddr_r_cry_1\);
    
    \rptr_gray[5]\ : SLE
      port map(D => \rptr_gray_1[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[5]_net_1\);
    
    fulli_0_a2_3 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[7]\, B => \wdiff_bus[8]\, C => 
        \wdiff_bus[9]\, D => \wdiff_bus[10]\, Y => \fulli_0_a2_3\);
    
    un1_memwaddr_r_s_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[12]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_11\, 
        S => un1_memwaddr_r_s_12_S, Y => OPEN, FCO => OPEN);
    
    \wptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[2]_net_1\, B => \wptr[3]_net_1\, Y => 
        \wptr_gray_1[2]_net_1\);
    
    \wptr[5]\ : SLE
      port map(D => \wptr_s[5]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => N_586, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr[5]_net_1\);
    
    rdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[5]_net_1\, B => 
        \rptr[5]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_4\, S => rdiff_bus(5), Y => OPEN, FCO => 
        \rdiff_bus_cry_5\);
    
    \wptr_bin_sync2[8]\ : SLE
      port map(D => \wptr_bin_sync[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[8]_net_1\);
    
    overflow_r_RNI5I9B : CFG1
      generic map(INIT => "01")

      port map(A => \RX_FIFO_OVERFLOW\, Y => RX_FIFO_OVERFLOW_i);
    
    \wptr[7]\ : SLE
      port map(D => \wptr_s[7]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => N_586, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr[7]_net_1\);
    
    un1_memwaddr_r_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_1\, 
        S => un1_memwaddr_r_cry_2_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_2\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \wptr_gray[1]\ : SLE
      port map(D => \wptr_gray_1[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[1]_net_1\);
    
    \rptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[9]_net_1\, B => \rptr[10]_net_1\, Y => 
        \rptr_gray_1[9]_net_1\);
    
    \rptr_bin_sync2[5]\ : SLE
      port map(D => \rptr_bin_sync[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[5]_net_1\);
    
    \rptr_bin_sync2[1]\ : SLE
      port map(D => \rptr_bin_sync[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[1]_net_1\);
    
    \memwaddr_r[10]\ : SLE
      port map(D => \memwaddr_r_2[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[10]\);
    
    wdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[7]_net_1\, B => 
        \rptr_bin_sync2[7]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_6\, S => \wdiff_bus[7]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_7\);
    
    \wptr_bin_sync2[0]\ : SLE
      port map(D => \wptr_bin_sync[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdiff_bus\);
    
    un1_memwaddr_r_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_7\, 
        S => un1_memwaddr_r_cry_8_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_8\);
    
    \wptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[0]_net_1\, S
         => \wptr_s[1]\, Y => OPEN, FCO => \wptr_cry[1]_net_1\);
    
    un1_memwaddr_r_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_3\, 
        S => un1_memwaddr_r_cry_4_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_4\);
    
    un1_memwaddr_r_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_2\, 
        S => un1_memwaddr_r_cry_3_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_3\);
    
    \memraddr_r[8]\ : SLE
      port map(D => \memraddr_r_2[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_283_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[8]\);
    
    \rptr[9]\ : SLE
      port map(D => \rptr_s[9]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => N_283_i, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[9]_net_1\);
    
    \wptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[6]_net_1\, B => \wptr[7]_net_1\, Y => 
        \wptr_gray_1[6]_net_1\);
    
    \wptr_gray[12]\ : SLE
      port map(D => \wptr_gray_1[12]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[12]_net_1\);
    
    \wptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[6]_net_1\, S
         => \wptr_s[7]\, Y => OPEN, FCO => \wptr_cry[7]_net_1\);
    
    \wptr_bin_sync2[2]\ : SLE
      port map(D => \wptr_bin_sync[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[2]_net_1\);
    
    fulli_0_1 : CFG4
      generic map(INIT => x"5557")

      port map(A => \fulli_0_a2_3\, B => N_567, C => 
        \wdiff_bus[5]\, D => \wdiff_bus[6]\, Y => \fulli_0_1\);
    
    \L1.un4_re_i_9\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \fifo_MEMRADDR[6]\, B => \fifo_MEMRADDR[5]\, 
        C => \fifo_MEMRADDR[0]\, D => un4_re_i_0, Y => un4_re_i_9);
    
    un1_memraddr_r_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_2\, 
        S => un1_memraddr_r_cry_3_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_3\);
    
    \rptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \rptr[0]_net_1\, Y => \rptr_s[0]\);
    
    un1_memraddr_r_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        un1_memraddr_r_s_1_275_FCO, S => un1_memraddr_r_cry_1_S, 
        Y => OPEN, FCO => \un1_memraddr_r_cry_1\);
    
    \rptr[4]\ : SLE
      port map(D => \rptr_s[4]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => N_283_i, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[4]_net_1\);
    
    \memwaddr_r_2[5]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_5_S, D => un4_we_i_9, Y => 
        \memwaddr_r_2[5]_net_1\);
    
    \wptr_gray[6]\ : SLE
      port map(D => \wptr_gray_1[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[6]_net_1\);
    
    \wptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[3]_net_1\, B => \wptr[4]_net_1\, Y => 
        \wptr_gray_1[3]_net_1\);
    
    \wptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[4]_net_1\, S
         => \wptr_s[5]\, Y => OPEN, FCO => \wptr_cry[5]_net_1\);
    
    un1_memraddr_r_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_8\, 
        S => un1_memraddr_r_cry_9_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_9\);
    
    \rptr_gray[4]\ : SLE
      port map(D => \rptr_gray_1[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[4]_net_1\);
    
    un1_memraddr_r_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_4\, 
        S => un1_memraddr_r_cry_5_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_5\);
    
    \wptr_bin_sync2[4]\ : SLE
      port map(D => bin_N_6_i_0, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr_bin_sync2[4]_net_1\);
    
    \wptr[3]\ : SLE
      port map(D => \wptr_s[3]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => N_586, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr[3]_net_1\);
    
    \L1.un4_we_i_9\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMWADDR[2]\, B => \fifo_MEMWADDR[1]\, 
        C => \fifo_MEMWADDR[0]\, D => un4_we_i_0, Y => un4_we_i_9);
    
    \memwaddr_r[6]\ : SLE
      port map(D => un1_memwaddr_r_cry_6_S, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[6]\);
    
    memwe_0_a2 : CFG2
      generic map(INIT => x"2")

      port map(A => N_586, B => \RX_FIFO_Full\, Y => \fifo_MEMWE\);
    
    \wptr[6]\ : SLE
      port map(D => \wptr_s[6]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => N_586, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr[6]_net_1\);
    
    \memwaddr_r[9]\ : SLE
      port map(D => \memwaddr_r_2[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[9]\);
    
    \memraddr_r[10]\ : SLE
      port map(D => \memraddr_r_2[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_283_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[10]\);
    
    \L1.un4_re_i_8\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMRADDR[12]\, B => \fifo_MEMRADDR[11]\, 
        C => \fifo_MEMRADDR[10]\, D => \fifo_MEMRADDR[9]\, Y => 
        un4_re_i_8);
    
    \memwaddr_r[3]\ : SLE
      port map(D => un1_memwaddr_r_cry_3_S, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[3]\);
    
    \rptr_gray_1[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[13]_net_1\, B => \rptr[12]_net_1\, Y
         => \rptr_gray_1[12]_net_1\);
    
    full_r : SLE
      port map(D => fulli, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_Full\);
    
    \rptr_bin_sync2[3]\ : SLE
      port map(D => \rptr_bin_sync[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[3]_net_1\);
    
    \rptr[2]\ : SLE
      port map(D => \rptr_s[2]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => N_283_i, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[2]_net_1\);
    
    \memraddr_r[3]\ : SLE
      port map(D => un1_memraddr_r_cry_3_S, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_283_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[3]\);
    
    \wptr_cry[0]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => wptr_cry_cy, S => 
        \wptr_s[0]\, Y => OPEN, FCO => \wptr_cry[0]_net_1\);
    
    \wptr[13]\ : SLE
      port map(D => \wptr_s[13]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_586, ALn => irx_fifo_rst_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \wptr[13]_net_1\);
    
    \rptr_bin_sync2[9]\ : SLE
      port map(D => \rptr_bin_sync[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[9]_net_1\);
    
    \wptr_bin_sync2[13]\ : SLE
      port map(D => \wptr_bin_sync[13]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[13]_net_1\);
    
    \rptr[11]\ : SLE
      port map(D => \rptr_s[11]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_283_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[11]_net_1\);
    
    \wptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[5]_net_1\, S
         => \wptr_s[6]\, Y => OPEN, FCO => \wptr_cry[6]_net_1\);
    
    \rptr_bin_sync2[11]\ : SLE
      port map(D => \rptr_bin_sync[11]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[11]_net_1\);
    
    \wptr_bin_sync2[5]\ : SLE
      port map(D => \wptr_bin_sync[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[5]_net_1\);
    
    \L1.un4_we_i_8\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMWADDR[8]\, B => \fifo_MEMWADDR[7]\, 
        C => \fifo_MEMWADDR[4]\, D => \fifo_MEMWADDR[3]\, Y => 
        un4_we_i_8);
    
    \wptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[7]_net_1\, S
         => \wptr_s[8]\, Y => OPEN, FCO => \wptr_cry[8]_net_1\);
    
    \wptr_bin_sync2[1]\ : SLE
      port map(D => \wptr_bin_sync[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[1]_net_1\);
    
    Wr_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_0
      port map(wptr_bin_sync(13) => \wptr_bin_sync[13]\, 
        wptr_bin_sync(12) => \wptr_bin_sync[12]\, 
        wptr_bin_sync(11) => \wptr_bin_sync[11]\, 
        wptr_bin_sync(10) => \wptr_bin_sync[10]\, 
        wptr_bin_sync(9) => \wptr_bin_sync[9]\, wptr_bin_sync(8)
         => \wptr_bin_sync[8]\, wptr_bin_sync(7) => 
        \wptr_bin_sync[7]\, wptr_bin_sync(6) => 
        \wptr_bin_sync[6]\, wptr_bin_sync(5) => 
        \wptr_bin_sync[5]\, wptr_bin_sync(4) => nc2, 
        wptr_bin_sync(3) => \wptr_bin_sync[3]\, wptr_bin_sync(2)
         => \wptr_bin_sync[2]\, wptr_bin_sync(1) => 
        \wptr_bin_sync[1]\, wptr_bin_sync(0) => 
        \wptr_bin_sync[0]\, wptr_gray_sync(12) => 
        \wptr_gray_sync[12]\, wptr_gray_sync(11) => 
        \wptr_gray_sync[11]\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\, bin_N_6_i => bin_N_6_i_0);
    
    \wptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[4]_net_1\, B => \wptr[5]_net_1\, Y => 
        \wptr_gray_1[4]_net_1\);
    
    \rptr_bin_sync2[13]\ : SLE
      port map(D => \rptr_bin_sync[13]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[13]_net_1\);
    
    \L1.un4_re_i_7\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMRADDR[8]\, B => \fifo_MEMRADDR[7]\, 
        C => \fifo_MEMRADDR[4]\, D => \fifo_MEMRADDR[3]\, Y => 
        un4_re_i_7);
    
    overflow_r : SLE
      port map(D => un1_we_p, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_OVERFLOW\);
    
    fulli_0 : CFG4
      generic map(INIT => x"BAAA")

      port map(A => \wdiff_bus[13]\, B => \fulli_0_1\, C => 
        \wdiff_bus[11]\, D => \wdiff_bus[12]\, Y => fulli);
    
    \memraddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMRADDR[0]\, Y => \fifo_MEMRADDR_i[0]\);
    
    \memraddr_r_2[8]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_8_S, D => un4_re_i_9, Y => 
        \memraddr_r_2[8]_net_1\);
    
    \rptr_gray[11]\ : SLE
      port map(D => \rptr_gray_1[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[10]\ : SLE
      port map(D => \wptr_bin_sync[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[10]_net_1\);
    
    \rptr[10]\ : SLE
      port map(D => \rptr_s[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_283_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[10]_net_1\);
    
    \wptr[9]\ : SLE
      port map(D => \wptr_s[9]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => N_586, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr[9]_net_1\);
    
    Wr_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1
      port map(wptr_gray(13) => \wptr_gray[13]_net_1\, 
        wptr_gray(12) => \wptr_gray[12]_net_1\, wptr_gray(11) => 
        \wptr_gray[11]_net_1\, wptr_gray(10) => 
        \wptr_gray[10]_net_1\, wptr_gray(9) => 
        \wptr_gray[9]_net_1\, wptr_gray(8) => 
        \wptr_gray[8]_net_1\, wptr_gray(7) => 
        \wptr_gray[7]_net_1\, wptr_gray(6) => 
        \wptr_gray[6]_net_1\, wptr_gray(5) => 
        \wptr_gray[5]_net_1\, wptr_gray(4) => 
        \wptr_gray[4]_net_1\, wptr_gray(3) => 
        \wptr_gray[3]_net_1\, wptr_gray(2) => 
        \wptr_gray[2]_net_1\, wptr_gray(1) => 
        \wptr_gray[1]_net_1\, wptr_gray(0) => 
        \wptr_gray[0]_net_1\, wptr_gray_sync(12) => 
        \wptr_gray_sync[12]\, wptr_gray_sync(11) => 
        \wptr_gray_sync[11]\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\, wptr_bin_sync_0 => 
        \wptr_bin_sync[13]\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, irx_fifo_rst_i => 
        irx_fifo_rst_i);
    
    un1_memwaddr_r_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_4\, 
        S => un1_memwaddr_r_cry_5_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_5\);
    
    \rptr_gray[0]\ : SLE
      port map(D => \rptr_gray_1[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[0]_net_1\);
    
    empty_r : SLE
      port map(D => empty_r_3, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => RX_FIFO_Empty);
    
    \memwaddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMWADDR[0]\, Y => \fifo_MEMWADDR_i[0]\);
    
    \memwaddr_r_2[12]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_s_12_S, D => un4_we_i_9, Y => 
        \memwaddr_r_2[12]_net_1\);
    
    \rptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[7]_net_1\, B => \rptr[8]_net_1\, Y => 
        \rptr_gray_1[7]_net_1\);
    
    un1_memraddr_r_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_1\, 
        S => un1_memraddr_r_cry_2_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_2\);
    
    wdiff_bus_cry_12 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[12]_net_1\, B => 
        \rptr_bin_sync2[12]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_11\, S => 
        \wdiff_bus[12]\, Y => OPEN, FCO => \wdiff_bus_cry_12\);
    
    \wptr[4]\ : SLE
      port map(D => \wptr_s[4]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => N_586, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr[4]_net_1\);
    
    un1_memraddr_r_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_7\, 
        S => un1_memraddr_r_cry_8_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_8\);
    
    \rptr_s[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[12]_net_1\, S
         => \rptr_s[13]_net_1\, Y => OPEN, FCO => OPEN);
    
    \memwaddr_r[8]\ : SLE
      port map(D => \memwaddr_r_2[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[8]\);
    
    \memwaddr_r[2]\ : SLE
      port map(D => un1_memwaddr_r_cry_2_S, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[2]\);
    
    \wptr_bin_sync2[11]\ : SLE
      port map(D => \wptr_bin_sync[11]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[11]_net_1\);
    
    \L1.un4_we_i_7\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \fifo_MEMWADDR[11]\, B => \fifo_MEMWADDR[10]\, 
        C => \fifo_MEMWADDR[9]\, D => \fifo_MEMWADDR[6]\, Y => 
        un4_we_i_7);
    
    \wptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[1]_net_1\, B => \wptr[2]_net_1\, Y => 
        \wptr_gray_1[1]_net_1\);
    
    underflow_r : SLE
      port map(D => un2_re_p, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RX_FIFO_UNDERRUN\);
    
    \memwaddr_r_2[11]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_11_S, D => un4_we_i_9, Y => 
        \memwaddr_r_2[11]_net_1\);
    
    \memraddr_r_2[12]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_s_12_S, D => un4_re_i_9, Y => 
        \memraddr_r_2[12]_net_1\);
    
    \wptr_gray[5]\ : SLE
      port map(D => \wptr_gray_1[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[5]_net_1\);
    
    \memraddr_r[7]\ : SLE
      port map(D => \memraddr_r_2[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_283_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[7]\);
    
    \L1.un1_we_p_0_a2\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_586, B => \RX_FIFO_Full\, Y => un1_we_p);
    
    un1_memraddr_r_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_5\, 
        S => un1_memraddr_r_cry_6_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_6\);
    
    \rptr_bin_sync2[10]\ : SLE
      port map(D => \rptr_bin_sync[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[10]_net_1\);
    
    wdiff_bus_s_13 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr_bin_sync2[13]_net_1\, C
         => \wptr[13]_net_1\, D => GND_net_1, FCI => 
        \wdiff_bus_cry_12\, S => \wdiff_bus[13]\, Y => OPEN, FCO
         => OPEN);
    
    wdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[10]_net_1\, B => 
        \rptr_bin_sync2[10]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_9\, S => \wdiff_bus[10]\, 
        Y => OPEN, FCO => \wdiff_bus_cry_10\);
    
    \memwaddr_r[11]\ : SLE
      port map(D => \memwaddr_r_2[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[11]\);
    
    \wptr_gray[8]\ : SLE
      port map(D => \wptr_gray_1[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[8]_net_1\);
    
    \memraddr_r_2[11]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_11_S, D => un4_re_i_9, Y => 
        \memraddr_r_2[11]_net_1\);
    
    un1_memraddr_r_s_1_275 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => un1_memraddr_r_s_1_275_FCO);
    
    un1_memraddr_r_s_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[12]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_11\, 
        S => un1_memraddr_r_s_12_S, Y => OPEN, FCO => OPEN);
    
    \wptr_gray[7]\ : SLE
      port map(D => \wptr_gray_1[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[7]_net_1\);
    
    \wptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[5]_net_1\, B => \wptr[6]_net_1\, Y => 
        \wptr_gray_1[5]_net_1\);
    
    \memwaddr_r[5]\ : SLE
      port map(D => \memwaddr_r_2[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[5]\);
    
    un1_memraddr_r_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_3\, 
        S => un1_memraddr_r_cry_4_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_4\);
    
    \rptr[8]\ : SLE
      port map(D => \rptr_s[8]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => N_283_i, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[8]_net_1\);
    
    Rd_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0
      port map(rptr_gray(13) => \rptr_gray[13]_net_1\, 
        rptr_gray(12) => \rptr_gray[12]_net_1\, rptr_gray(11) => 
        \rptr_gray[11]_net_1\, rptr_gray(10) => 
        \rptr_gray[10]_net_1\, rptr_gray(9) => 
        \rptr_gray[9]_net_1\, rptr_gray(8) => 
        \rptr_gray[8]_net_1\, rptr_gray(7) => 
        \rptr_gray[7]_net_1\, rptr_gray(6) => 
        \rptr_gray[6]_net_1\, rptr_gray(5) => 
        \rptr_gray[5]_net_1\, rptr_gray(4) => 
        \rptr_gray[4]_net_1\, rptr_gray(3) => 
        \rptr_gray[3]_net_1\, rptr_gray(2) => 
        \rptr_gray[2]_net_1\, rptr_gray(1) => 
        \rptr_gray[1]_net_1\, rptr_gray(0) => 
        \rptr_gray[0]_net_1\, rptr_gray_sync(12) => 
        \rptr_gray_sync[12]\, rptr_gray_sync(11) => 
        \rptr_gray_sync[11]\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\, rptr_bin_sync_0 => 
        \rptr_bin_sync[13]\, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, irx_fifo_rst_i => irx_fifo_rst_i);
    
    \rptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[3]_net_1\, S
         => \rptr_s[4]\, Y => OPEN, FCO => \rptr_cry[4]_net_1\);
    
    wdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[2]_net_1\, B => 
        \rptr_bin_sync2[2]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_1\, S => \wdiff_bus[2]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_2\);
    
    \rptr_gray[2]\ : SLE
      port map(D => \rptr_gray_1[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[2]_net_1\);
    
    \wptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[8]_net_1\, S
         => \wptr_s[9]\, Y => OPEN, FCO => \wptr_cry[9]_net_1\);
    
    \wptr_bin_sync2[3]\ : SLE
      port map(D => \wptr_bin_sync[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[3]_net_1\);
    
    \rptr[12]\ : SLE
      port map(D => \rptr_s[12]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_283_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[12]_net_1\);
    
    \wptr[2]\ : SLE
      port map(D => \wptr_s[2]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => N_586, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr[2]_net_1\);
    
    \rptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[1]_net_1\, S
         => \rptr_s[2]\, Y => OPEN, FCO => \rptr_cry[2]_net_1\);
    
    rdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[9]_net_1\, B => 
        \rptr[9]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_8\, S => rdiff_bus(9), Y => OPEN, FCO => 
        \rdiff_bus_cry_9\);
    
    \memwaddr_r[0]\ : SLE
      port map(D => \fifo_MEMWADDR_i[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[0]\);
    
    \wptr_gray[2]\ : SLE
      port map(D => \wptr_gray_1[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[2]_net_1\);
    
    \wptr_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[11]_net_1\, S
         => \wptr_s[12]\, Y => OPEN, FCO => \wptr_cry[12]_net_1\);
    
    \memwaddr_r_2[7]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_7_S, D => un4_we_i_9, Y => 
        \memwaddr_r_2[7]_net_1\);
    
    wdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[4]_net_1\, B => 
        \rptr_bin_sync2[4]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_3\, S => \wdiff_bus[4]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_4\);
    
    un1_memraddr_r_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_6\, 
        S => un1_memraddr_r_cry_7_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_7\);
    
    \wptr_s[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[12]_net_1\, S
         => \wptr_s[13]_net_1\, Y => OPEN, FCO => OPEN);
    
    \wptr_gray[11]\ : SLE
      port map(D => \wptr_gray_1[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[9]\ : SLE
      port map(D => \wptr_bin_sync[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[9]_net_1\);
    
    \wptr_cry_cy[0]\ : ARI1
      generic map(INIT => x"45500")

      port map(A => VCC_net_1, B => \RX_FIFO_Full\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => wptr_cry_cy);
    
    \rptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[6]_net_1\, B => \rptr[7]_net_1\, Y => 
        \rptr_gray_1[6]_net_1\);
    
    \wptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[10]_net_1\, B => \wptr[11]_net_1\, Y
         => \wptr_gray_1[10]_net_1\);
    
    wdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[6]_net_1\, B => 
        \rptr_bin_sync2[6]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_5\, S => \wdiff_bus[6]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_6\);
    
    \rptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[2]_net_1\, S
         => \rptr_s[3]\, Y => OPEN, FCO => \rptr_cry[3]_net_1\);
    
    \memraddr_r[4]\ : SLE
      port map(D => un1_memraddr_r_cry_4_S, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_283_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[4]\);
    
    \rptr[13]\ : SLE
      port map(D => \rptr_s[13]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_283_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[13]_net_1\);
    
    \wptr_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[10]_net_1\, S
         => \wptr_s[11]\, Y => OPEN, FCO => \wptr_cry[11]_net_1\);
    
    \memwaddr_r_2[8]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_8_S, D => un4_we_i_9, Y => 
        \memwaddr_r_2[8]_net_1\);
    
    \memwaddr_r[12]\ : SLE
      port map(D => \memwaddr_r_2[12]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[12]\);
    
    \L1.un4_re_i_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \fifo_MEMRADDR[1]\, B => \fifo_MEMRADDR[2]\, 
        Y => un4_re_i_0);
    
    \rptr_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[11]_net_1\, S
         => \rptr_s[12]\, Y => OPEN, FCO => \rptr_cry[12]_net_1\);
    
    \memraddr_r[11]\ : SLE
      port map(D => \memraddr_r_2[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_283_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[11]\);
    
    rdiff_bus_cry_12 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[12]_net_1\, B => 
        \rptr[12]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_11\, S => rdiff_bus(12), Y => OPEN, FCO
         => \rdiff_bus_cry_12\);
    
    \memraddr_r[5]\ : SLE
      port map(D => \memraddr_r_2[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_283_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[5]\);
    
    \rptr_gray[6]\ : SLE
      port map(D => \rptr_gray_1[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[6]_net_1\);
    
    \memraddr_r[9]\ : SLE
      port map(D => \memraddr_r_2[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_283_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[9]\);
    
    \rptr[0]\ : SLE
      port map(D => \rptr_s[0]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => N_283_i, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[0]_net_1\);
    
    \wptr[10]\ : SLE
      port map(D => \wptr_s[10]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => N_586, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr[10]_net_1\);
    
    \L1.un4_we_i_0\ : CFG2
      generic map(INIT => x"4")

      port map(A => \fifo_MEMWADDR[5]\, B => \fifo_MEMWADDR[12]\, 
        Y => un4_we_i_0);
    
    wdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[1]_net_1\, B => 
        \rptr_bin_sync2[1]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_0\, S => \wdiff_bus[1]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_1\);
    
    rdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[2]_net_1\, B => 
        \rptr[2]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_1\, S => rdiff_bus(2), Y => OPEN, FCO => 
        \rdiff_bus_cry_2\);
    
    \wptr_gray[9]\ : SLE
      port map(D => \wptr_gray_1[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[9]_net_1\);
    
    \rptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[4]_net_1\, B => \rptr[5]_net_1\, Y => 
        \rptr_gray_1[4]_net_1\);
    
    fulli_0_a2_0_2 : CFG3
      generic map(INIT => x"20")

      port map(A => \wdiff_bus[4]\, B => wdiff_bus_cry_0_Y_0, C
         => \wdiff_bus[1]\, Y => \fulli_0_a2_0_2\);
    
    \wptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[8]_net_1\, B => \wptr[9]_net_1\, Y => 
        \wptr_gray_1[8]_net_1\);
    
    Rd_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv
      port map(rptr_bin_sync(13) => \rptr_bin_sync[13]\, 
        rptr_bin_sync(12) => \rptr_bin_sync[12]\, 
        rptr_bin_sync(11) => \rptr_bin_sync[11]\, 
        rptr_bin_sync(10) => \rptr_bin_sync[10]\, 
        rptr_bin_sync(9) => \rptr_bin_sync[9]\, rptr_bin_sync(8)
         => \rptr_bin_sync[8]\, rptr_bin_sync(7) => 
        \rptr_bin_sync[7]\, rptr_bin_sync(6) => 
        \rptr_bin_sync[6]\, rptr_bin_sync(5) => 
        \rptr_bin_sync[5]\, rptr_bin_sync(4) => nc1, 
        rptr_bin_sync(3) => \rptr_bin_sync[3]\, rptr_bin_sync(2)
         => \rptr_bin_sync[2]\, rptr_bin_sync(1) => 
        \rptr_bin_sync[1]\, rptr_bin_sync(0) => 
        \rptr_bin_sync[0]\, rptr_gray_sync(12) => 
        \rptr_gray_sync[12]\, rptr_gray_sync(11) => 
        \rptr_gray_sync[11]\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\, bin_N_6_i => bin_N_6_i);
    
    \rptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => rptr_s_266_FCO, S => 
        \rptr_s[1]\, Y => OPEN, FCO => \rptr_cry[1]_net_1\);
    
    \rptr_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[10]_net_1\, S
         => \rptr_s[11]\, Y => OPEN, FCO => \rptr_cry[11]_net_1\);
    
    rdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[3]_net_1\, B => 
        \rptr[3]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_2\, S => rdiff_bus(3), Y => OPEN, FCO => 
        \rdiff_bus_cry_3\);
    
    rdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[10]_net_1\, B => 
        \rptr[10]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_9\, S => rdiff_bus(10), Y => OPEN, FCO => 
        \rdiff_bus_cry_10\);
    
    un1_memwaddr_r_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[11]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_10\, 
        S => un1_memwaddr_r_cry_11_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_11\);
    
    \memraddr_r[6]\ : SLE
      port map(D => un1_memraddr_r_cry_6_S, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_283_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[6]\);
    
    \rptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[6]_net_1\, S
         => \rptr_s[7]\, Y => OPEN, FCO => \rptr_cry[7]_net_1\);
    
    rdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rdiff_bus\, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => rdiff_bus_cry_0_Y_0, FCO => \rdiff_bus_cry_0\);
    
    \memraddr_r[2]\ : SLE
      port map(D => un1_memraddr_r_cry_2_S, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_283_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[2]\);
    
    \wptr[8]\ : SLE
      port map(D => \wptr_s[8]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => N_586, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr[8]_net_1\);
    
    wdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[3]_net_1\, B => 
        \rptr_bin_sync2[3]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_2\, S => \wdiff_bus[3]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_3\);
    
    rdiff_bus_s_13 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr[13]_net_1\, C => 
        \wptr_bin_sync2[13]_net_1\, D => GND_net_1, FCI => 
        \rdiff_bus_cry_12\, S => rdiff_bus(13), Y => OPEN, FCO
         => OPEN);
    
    \memraddr_r[12]\ : SLE
      port map(D => \memraddr_r_2[12]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_283_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[12]\);
    
    \wptr_gray_1[11]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[11]_net_1\, B => \wptr[12]_net_1\, Y
         => \wptr_gray_1[11]_net_1\);
    
    \rptr_gray[7]\ : SLE
      port map(D => \rptr_gray_1[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[7]_net_1\);
    
    \wptr_gray[0]\ : SLE
      port map(D => \wptr_gray_1[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[0]_net_1\);
    
    \rptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[0]_net_1\, B => \rptr[1]_net_1\, Y => 
        \rptr_gray_1[0]_net_1\);
    
    un1_memwaddr_r_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_9\, 
        S => un1_memwaddr_r_cry_10_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_10\);
    
    \rptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[8]_net_1\, B => \rptr[9]_net_1\, Y => 
        \rptr_gray_1[8]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO is

    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          rdiff_bus                 : out   std_logic_vector(13 downto 1);
          RDATA_int                 : out   std_logic_vector(7 downto 0);
          RDATA_r                   : out   std_logic_vector(7 downto 0);
          RX_FIFO_UNDERRUN          : out   std_logic;
          RX_FIFO_UNDERRUN_i        : out   std_logic;
          RX_FIFO_OVERFLOW          : out   std_logic;
          RX_FIFO_OVERFLOW_i        : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          RX_FIFO_Empty             : out   std_logic;
          empty_r_3                 : in    std_logic;
          RX_FIFO_Full              : out   std_logic;
          un2_re_p                  : in    std_logic;
          rdiff_bus_cry_0_Y_0       : out   std_logic;
          iRX_FIFO_wr_en            : in    std_logic;
          sampler_clk1x_en          : in    std_logic;
          RX_InProcess_d1           : in    std_logic;
          tx_col_detect_en          : in    std_logic;
          N_357                     : out   std_logic;
          re_pulse_d1               : out   std_logic;
          RX_FIFO_rd_en             : in    std_logic;
          RE_d1                     : out   std_logic;
          N_283_i                   : in    std_logic;
          N_314_i_i                 : in    std_logic;
          REN_d1                    : out   std_logic;
          iRX_FIFO_rd_en_RNIJFNA_0  : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper
    port( fifo_MEMRADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          N_283_i                   : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          fifo_MEMWE                : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async
    port( rdiff_bus                 : out   std_logic_vector(13 downto 1);
          fifo_MEMRADDR             : out   std_logic_vector(12 downto 0);
          fifo_MEMWADDR             : out   std_logic_vector(12 downto 0);
          tx_col_detect_en          : in    std_logic := 'U';
          RX_InProcess_d1           : in    std_logic := 'U';
          sampler_clk1x_en          : in    std_logic := 'U';
          iRX_FIFO_wr_en            : in    std_logic := 'U';
          rdiff_bus_cry_0_Y_0       : out   std_logic;
          un2_re_p                  : in    std_logic := 'U';
          RX_FIFO_Full              : out   std_logic;
          empty_r_3                 : in    std_logic := 'U';
          RX_FIFO_Empty             : out   std_logic;
          N_283_i                   : in    std_logic := 'U';
          fifo_MEMWE                : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U';
          RX_FIFO_OVERFLOW_i        : out   std_logic;
          RX_FIFO_OVERFLOW          : out   std_logic;
          RX_FIFO_UNDERRUN_i        : out   std_logic;
          RX_FIFO_UNDERRUN          : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \RDATA_int[0]\, GND_net_1, \RDATA_int[1]\, 
        \RDATA_int[2]\, \RDATA_int[3]\, \RDATA_int[4]\, 
        \RDATA_int[5]\, \RDATA_int[6]\, \RDATA_int[7]\, 
        \RDATA_r[8]_net_1\, \RDATA_int[8]\, \re_set\, 
        REN_d1_net_1, RE_d1_net_1, re_pulse_d1_net_1, \re_pulse\, 
        \fifo_MEMRADDR[0]\, \fifo_MEMRADDR[1]\, 
        \fifo_MEMRADDR[2]\, \fifo_MEMRADDR[3]\, 
        \fifo_MEMRADDR[4]\, \fifo_MEMRADDR[5]\, 
        \fifo_MEMRADDR[6]\, \fifo_MEMRADDR[7]\, 
        \fifo_MEMRADDR[8]\, \fifo_MEMRADDR[9]\, 
        \fifo_MEMRADDR[10]\, \fifo_MEMRADDR[11]\, 
        \fifo_MEMRADDR[12]\, \fifo_MEMWADDR[0]\, 
        \fifo_MEMWADDR[1]\, \fifo_MEMWADDR[2]\, 
        \fifo_MEMWADDR[3]\, \fifo_MEMWADDR[4]\, 
        \fifo_MEMWADDR[5]\, \fifo_MEMWADDR[6]\, 
        \fifo_MEMWADDR[7]\, \fifo_MEMWADDR[8]\, 
        \fifo_MEMWADDR[9]\, \fifo_MEMWADDR[10]\, 
        \fifo_MEMWADDR[11]\, \fifo_MEMWADDR[12]\, fifo_MEMWE
         : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async(DEF_ARCH);
begin 

    RDATA_int(7) <= \RDATA_int[7]\;
    RDATA_int(6) <= \RDATA_int[6]\;
    RDATA_int(5) <= \RDATA_int[5]\;
    RDATA_int(4) <= \RDATA_int[4]\;
    RDATA_int(3) <= \RDATA_int[3]\;
    RDATA_int(2) <= \RDATA_int[2]\;
    RDATA_int(1) <= \RDATA_int[1]\;
    RDATA_int(0) <= \RDATA_int[0]\;
    re_pulse_d1 <= re_pulse_d1_net_1;
    RE_d1 <= RE_d1_net_1;
    REN_d1 <= REN_d1_net_1;

    re_pulse : CFG2
      generic map(INIT => x"E")

      port map(A => iRX_FIFO_rd_en_RNIJFNA_0, B => \re_set\, Y
         => \re_pulse\);
    
    \RDATA_r[3]\ : SLE
      port map(D => \RDATA_int[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => iRX_FIFO_rd_en_RNIJFNA_0, 
        ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => RDATA_r(3));
    
    \re_pulse_d1\ : SLE
      port map(D => \re_pulse\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => re_pulse_d1_net_1);
    
    \RDATA_r[5]\ : SLE
      port map(D => \RDATA_int[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => iRX_FIFO_rd_en_RNIJFNA_0, 
        ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => RDATA_r(5));
    
    \RDATA_r[8]\ : SLE
      port map(D => \RDATA_int[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => iRX_FIFO_rd_en_RNIJFNA_0, 
        ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[8]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \RW1.UI_ram_wrapper_1\ : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper
      port map(fifo_MEMRADDR(12) => \fifo_MEMRADDR[12]\, 
        fifo_MEMRADDR(11) => \fifo_MEMRADDR[11]\, 
        fifo_MEMRADDR(10) => \fifo_MEMRADDR[10]\, 
        fifo_MEMRADDR(9) => \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8)
         => \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, fifo_MEMWADDR(12) => 
        \fifo_MEMWADDR[12]\, fifo_MEMWADDR(11) => 
        \fifo_MEMWADDR[11]\, fifo_MEMWADDR(10) => 
        \fifo_MEMWADDR[10]\, fifo_MEMWADDR(9) => 
        \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8) => 
        \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, RDATA_int(8) => \RDATA_int[8]\, 
        RDATA_int(7) => \RDATA_int[7]\, RDATA_int(6) => 
        \RDATA_int[6]\, RDATA_int(5) => \RDATA_int[5]\, 
        RDATA_int(4) => \RDATA_int[4]\, RDATA_int(3) => 
        \RDATA_int[3]\, RDATA_int(2) => \RDATA_int[2]\, 
        RDATA_int(1) => \RDATA_int[1]\, RDATA_int(0) => 
        \RDATA_int[0]\, RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, N_283_i => N_283_i, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, fifo_MEMWE
         => fifo_MEMWE);
    
    \RDATA_r[0]\ : SLE
      port map(D => \RDATA_int[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => iRX_FIFO_rd_en_RNIJFNA_0, 
        ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => RDATA_r(0));
    
    \RDATA_r[2]\ : SLE
      port map(D => \RDATA_int[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => iRX_FIFO_rd_en_RNIJFNA_0, 
        ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => RDATA_r(2));
    
    \RDATA_r[6]\ : SLE
      port map(D => \RDATA_int[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => iRX_FIFO_rd_en_RNIJFNA_0, 
        ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => RDATA_r(6));
    
    \L31.U_corefifo_async\ : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async
      port map(rdiff_bus(13) => rdiff_bus(13), rdiff_bus(12) => 
        rdiff_bus(12), rdiff_bus(11) => rdiff_bus(11), 
        rdiff_bus(10) => rdiff_bus(10), rdiff_bus(9) => 
        rdiff_bus(9), rdiff_bus(8) => rdiff_bus(8), rdiff_bus(7)
         => rdiff_bus(7), rdiff_bus(6) => rdiff_bus(6), 
        rdiff_bus(5) => rdiff_bus(5), rdiff_bus(4) => 
        rdiff_bus(4), rdiff_bus(3) => rdiff_bus(3), rdiff_bus(2)
         => rdiff_bus(2), rdiff_bus(1) => rdiff_bus(1), 
        fifo_MEMRADDR(12) => \fifo_MEMRADDR[12]\, 
        fifo_MEMRADDR(11) => \fifo_MEMRADDR[11]\, 
        fifo_MEMRADDR(10) => \fifo_MEMRADDR[10]\, 
        fifo_MEMRADDR(9) => \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8)
         => \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, fifo_MEMWADDR(12) => 
        \fifo_MEMWADDR[12]\, fifo_MEMWADDR(11) => 
        \fifo_MEMWADDR[11]\, fifo_MEMWADDR(10) => 
        \fifo_MEMWADDR[10]\, fifo_MEMWADDR(9) => 
        \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8) => 
        \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, tx_col_detect_en => tx_col_detect_en, 
        RX_InProcess_d1 => RX_InProcess_d1, sampler_clk1x_en => 
        sampler_clk1x_en, iRX_FIFO_wr_en => iRX_FIFO_wr_en, 
        rdiff_bus_cry_0_Y_0 => rdiff_bus_cry_0_Y_0, un2_re_p => 
        un2_re_p, RX_FIFO_Full => RX_FIFO_Full, empty_r_3 => 
        empty_r_3, RX_FIFO_Empty => RX_FIFO_Empty, N_283_i => 
        N_283_i, fifo_MEMWE => fifo_MEMWE, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        irx_fifo_rst_i => irx_fifo_rst_i, RX_FIFO_OVERFLOW_i => 
        RX_FIFO_OVERFLOW_i, RX_FIFO_OVERFLOW => RX_FIFO_OVERFLOW, 
        RX_FIFO_UNDERRUN_i => RX_FIFO_UNDERRUN_i, 
        RX_FIFO_UNDERRUN => RX_FIFO_UNDERRUN);
    
    re_set : SLE
      port map(D => REN_d1_net_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_314_i_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \re_set\);
    
    \Q_i_m2[8]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => re_pulse_d1_net_1, B => \RDATA_r[8]_net_1\, C
         => \RDATA_int[8]\, D => RE_d1_net_1, Y => N_357);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \RE_d1\ : SLE
      port map(D => RX_FIFO_rd_en, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RE_d1_net_1);
    
    \RDATA_r[7]\ : SLE
      port map(D => \RDATA_int[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => iRX_FIFO_rd_en_RNIJFNA_0, 
        ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => RDATA_r(7));
    
    \RDATA_r[4]\ : SLE
      port map(D => \RDATA_int[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => iRX_FIFO_rd_en_RNIJFNA_0, 
        ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => RDATA_r(4));
    
    \REN_d1\ : SLE
      port map(D => N_283_i, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => REN_d1_net_1);
    
    \RDATA_r[1]\ : SLE
      port map(D => \RDATA_int[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => iRX_FIFO_rd_en_RNIJFNA_0, 
        ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => RDATA_r(1));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9 is

    port( RDATA_r                   : out   std_logic_vector(7 downto 0);
          RDATA_int                 : out   std_logic_vector(7 downto 0);
          rdiff_bus                 : out   std_logic_vector(13 downto 1);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          irx_fifo_rst_i            : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          iRX_FIFO_rd_en_RNIJFNA_0  : in    std_logic;
          REN_d1                    : out   std_logic;
          N_314_i_i                 : in    std_logic;
          N_283_i                   : in    std_logic;
          RE_d1                     : out   std_logic;
          RX_FIFO_rd_en             : in    std_logic;
          re_pulse_d1               : out   std_logic;
          N_357                     : out   std_logic;
          tx_col_detect_en          : in    std_logic;
          RX_InProcess_d1           : in    std_logic;
          sampler_clk1x_en          : in    std_logic;
          iRX_FIFO_wr_en            : in    std_logic;
          rdiff_bus_cry_0_Y_0       : out   std_logic;
          un2_re_p                  : in    std_logic;
          RX_FIFO_Full              : out   std_logic;
          empty_r_3                 : in    std_logic;
          RX_FIFO_Empty             : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          RX_FIFO_OVERFLOW_i        : out   std_logic;
          RX_FIFO_OVERFLOW          : out   std_logic;
          RX_FIFO_UNDERRUN_i        : out   std_logic;
          RX_FIFO_UNDERRUN          : out   std_logic
        );

end FIFO_8Kx9;

architecture DEF_ARCH of FIFO_8Kx9 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO
    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          rdiff_bus                 : out   std_logic_vector(13 downto 1);
          RDATA_int                 : out   std_logic_vector(7 downto 0);
          RDATA_r                   : out   std_logic_vector(7 downto 0);
          RX_FIFO_UNDERRUN          : out   std_logic;
          RX_FIFO_UNDERRUN_i        : out   std_logic;
          RX_FIFO_OVERFLOW          : out   std_logic;
          RX_FIFO_OVERFLOW_i        : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          RX_FIFO_Empty             : out   std_logic;
          empty_r_3                 : in    std_logic := 'U';
          RX_FIFO_Full              : out   std_logic;
          un2_re_p                  : in    std_logic := 'U';
          rdiff_bus_cry_0_Y_0       : out   std_logic;
          iRX_FIFO_wr_en            : in    std_logic := 'U';
          sampler_clk1x_en          : in    std_logic := 'U';
          RX_InProcess_d1           : in    std_logic := 'U';
          tx_col_detect_en          : in    std_logic := 'U';
          N_357                     : out   std_logic;
          re_pulse_d1               : out   std_logic;
          RX_FIFO_rd_en             : in    std_logic := 'U';
          RE_d1                     : out   std_logic;
          N_283_i                   : in    std_logic := 'U';
          N_314_i_i                 : in    std_logic := 'U';
          REN_d1                    : out   std_logic;
          iRX_FIFO_rd_en_RNIJFNA_0  : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    FIFO_8Kx9_0 : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO
      port map(RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), rdiff_bus(13)
         => rdiff_bus(13), rdiff_bus(12) => rdiff_bus(12), 
        rdiff_bus(11) => rdiff_bus(11), rdiff_bus(10) => 
        rdiff_bus(10), rdiff_bus(9) => rdiff_bus(9), rdiff_bus(8)
         => rdiff_bus(8), rdiff_bus(7) => rdiff_bus(7), 
        rdiff_bus(6) => rdiff_bus(6), rdiff_bus(5) => 
        rdiff_bus(5), rdiff_bus(4) => rdiff_bus(4), rdiff_bus(3)
         => rdiff_bus(3), rdiff_bus(2) => rdiff_bus(2), 
        rdiff_bus(1) => rdiff_bus(1), RDATA_int(7) => 
        RDATA_int(7), RDATA_int(6) => RDATA_int(6), RDATA_int(5)
         => RDATA_int(5), RDATA_int(4) => RDATA_int(4), 
        RDATA_int(3) => RDATA_int(3), RDATA_int(2) => 
        RDATA_int(2), RDATA_int(1) => RDATA_int(1), RDATA_int(0)
         => RDATA_int(0), RDATA_r(7) => RDATA_r(7), RDATA_r(6)
         => RDATA_r(6), RDATA_r(5) => RDATA_r(5), RDATA_r(4) => 
        RDATA_r(4), RDATA_r(3) => RDATA_r(3), RDATA_r(2) => 
        RDATA_r(2), RDATA_r(1) => RDATA_r(1), RDATA_r(0) => 
        RDATA_r(0), RX_FIFO_UNDERRUN => RX_FIFO_UNDERRUN, 
        RX_FIFO_UNDERRUN_i => RX_FIFO_UNDERRUN_i, 
        RX_FIFO_OVERFLOW => RX_FIFO_OVERFLOW, RX_FIFO_OVERFLOW_i
         => RX_FIFO_OVERFLOW_i, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, RX_FIFO_Empty => RX_FIFO_Empty, 
        empty_r_3 => empty_r_3, RX_FIFO_Full => RX_FIFO_Full, 
        un2_re_p => un2_re_p, rdiff_bus_cry_0_Y_0 => 
        rdiff_bus_cry_0_Y_0, iRX_FIFO_wr_en => iRX_FIFO_wr_en, 
        sampler_clk1x_en => sampler_clk1x_en, RX_InProcess_d1 => 
        RX_InProcess_d1, tx_col_detect_en => tx_col_detect_en, 
        N_357 => N_357, re_pulse_d1 => re_pulse_d1, RX_FIFO_rd_en
         => RX_FIFO_rd_en, RE_d1 => RE_d1, N_283_i => N_283_i, 
        N_314_i_i => N_314_i_i, REN_d1 => REN_d1, 
        iRX_FIFO_rd_en_RNIJFNA_0 => iRX_FIFO_rd_en_RNIJFNA_0, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        irx_fifo_rst_i => irx_fifo_rst_i);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top is

    port( fifo_MEMWADDR                : in    std_logic_vector(10 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          fifo_MEMRADDR                : in    std_logic_vector(10 downto 0);
          RDATA_int                    : out   std_logic_vector(7 downto 0);
          fifo_MEMWE                   : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic;
          fifo_MEMRE                   : in    std_logic;
          BIT_CLK                      : in    std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top;

architecture DEF_ARCH of FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component RAM1K18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_CLK         : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ARST_N      : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          A_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_CLK         : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ARST_N      : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          B_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_WMODE       : in    std_logic := 'U';
          B_EN          : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_WMODE       : in    std_logic := 'U';
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;
    signal nc24, nc1, nc8, nc13, nc16, nc19, nc25, nc20, nc27, 
        nc9, nc22, nc28, nc14, nc5, nc21, nc15, nc3, nc10, nc7, 
        nc17, nc4, nc12, nc2, nc23, nc18, nc26, nc6, nc11
         : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top_R0C0 : RAM1K18
      port map(A_DOUT(17) => nc24, A_DOUT(16) => nc1, A_DOUT(15)
         => nc8, A_DOUT(14) => nc13, A_DOUT(13) => nc16, 
        A_DOUT(12) => nc19, A_DOUT(11) => nc25, A_DOUT(10) => 
        nc20, A_DOUT(9) => nc27, A_DOUT(8) => nc9, A_DOUT(7) => 
        RDATA_int(7), A_DOUT(6) => RDATA_int(6), A_DOUT(5) => 
        RDATA_int(5), A_DOUT(4) => RDATA_int(4), A_DOUT(3) => 
        RDATA_int(3), A_DOUT(2) => RDATA_int(2), A_DOUT(1) => 
        RDATA_int(1), A_DOUT(0) => RDATA_int(0), B_DOUT(17) => 
        nc22, B_DOUT(16) => nc28, B_DOUT(15) => nc14, B_DOUT(14)
         => nc5, B_DOUT(13) => nc21, B_DOUT(12) => nc15, 
        B_DOUT(11) => nc3, B_DOUT(10) => nc10, B_DOUT(9) => nc7, 
        B_DOUT(8) => nc17, B_DOUT(7) => nc4, B_DOUT(6) => nc12, 
        B_DOUT(5) => nc2, B_DOUT(4) => nc23, B_DOUT(3) => nc18, 
        B_DOUT(2) => nc26, B_DOUT(1) => nc6, B_DOUT(0) => nc11, 
        BUSY => OPEN, A_CLK => BIT_CLK, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(10), A_ADDR(12) => fifo_MEMRADDR(9), 
        A_ADDR(11) => fifo_MEMRADDR(8), A_ADDR(10) => 
        fifo_MEMRADDR(7), A_ADDR(9) => fifo_MEMRADDR(6), 
        A_ADDR(8) => fifo_MEMRADDR(5), A_ADDR(7) => 
        fifo_MEMRADDR(4), A_ADDR(6) => fifo_MEMRADDR(3), 
        A_ADDR(5) => fifo_MEMRADDR(2), A_ADDR(4) => 
        fifo_MEMRADDR(1), A_ADDR(3) => fifo_MEMRADDR(0), 
        A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, A_ADDR(0)
         => GND_net_1, A_WEN(1) => GND_net_1, A_WEN(0) => 
        GND_net_1, B_CLK => m2s010_som_sb_0_CCC_71MHz, B_DOUT_CLK
         => VCC_net_1, B_ARST_N => VCC_net_1, B_DOUT_EN => 
        VCC_net_1, B_BLK(2) => fifo_MEMWE, B_BLK(1) => VCC_net_1, 
        B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => GND_net_1, 
        B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => GND_net_1, 
        B_DIN(16) => GND_net_1, B_DIN(15) => GND_net_1, B_DIN(14)
         => GND_net_1, B_DIN(13) => GND_net_1, B_DIN(12) => 
        GND_net_1, B_DIN(11) => GND_net_1, B_DIN(10) => GND_net_1, 
        B_DIN(9) => GND_net_1, B_DIN(8) => GND_net_1, B_DIN(7)
         => CoreAPB3_0_APBmslave0_PWDATA(7), B_DIN(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), B_DIN(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), B_DIN(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), B_DIN(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), B_DIN(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), B_DIN(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), B_DIN(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), B_ADDR(13) => 
        fifo_MEMWADDR(10), B_ADDR(12) => fifo_MEMWADDR(9), 
        B_ADDR(11) => fifo_MEMWADDR(8), B_ADDR(10) => 
        fifo_MEMWADDR(7), B_ADDR(9) => fifo_MEMWADDR(6), 
        B_ADDR(8) => fifo_MEMWADDR(5), B_ADDR(7) => 
        fifo_MEMWADDR(4), B_ADDR(6) => fifo_MEMWADDR(3), 
        B_ADDR(5) => fifo_MEMWADDR(2), B_ADDR(4) => 
        fifo_MEMWADDR(1), B_ADDR(3) => fifo_MEMWADDR(0), 
        B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, B_ADDR(0)
         => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0) => 
        VCC_net_1, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper is

    port( RDATA_int                    : out   std_logic_vector(7 downto 0);
          fifo_MEMRADDR                : in    std_logic_vector(10 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          fifo_MEMWADDR                : in    std_logic_vector(10 downto 0);
          BIT_CLK                      : in    std_logic;
          fifo_MEMRE                   : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic;
          fifo_MEMWE                   : in    std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper;

architecture DEF_ARCH of FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top
    port( fifo_MEMWADDR                : in    std_logic_vector(10 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          fifo_MEMRADDR                : in    std_logic_vector(10 downto 0) := (others => 'U');
          RDATA_int                    : out   std_logic_vector(7 downto 0);
          fifo_MEMWE                   : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic := 'U';
          fifo_MEMRE                   : in    std_logic := 'U';
          BIT_CLK                      : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top
	Use entity work.FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    L1_asyncnonpipe : FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top
      port map(fifo_MEMWADDR(10) => fifo_MEMWADDR(10), 
        fifo_MEMWADDR(9) => fifo_MEMWADDR(9), fifo_MEMWADDR(8)
         => fifo_MEMWADDR(8), fifo_MEMWADDR(7) => 
        fifo_MEMWADDR(7), fifo_MEMWADDR(6) => fifo_MEMWADDR(6), 
        fifo_MEMWADDR(5) => fifo_MEMWADDR(5), fifo_MEMWADDR(4)
         => fifo_MEMWADDR(4), fifo_MEMWADDR(3) => 
        fifo_MEMWADDR(3), fifo_MEMWADDR(2) => fifo_MEMWADDR(2), 
        fifo_MEMWADDR(1) => fifo_MEMWADDR(1), fifo_MEMWADDR(0)
         => fifo_MEMWADDR(0), CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), fifo_MEMRADDR(10) => 
        fifo_MEMRADDR(10), fifo_MEMRADDR(9) => fifo_MEMRADDR(9), 
        fifo_MEMRADDR(8) => fifo_MEMRADDR(8), fifo_MEMRADDR(7)
         => fifo_MEMRADDR(7), fifo_MEMRADDR(6) => 
        fifo_MEMRADDR(6), fifo_MEMRADDR(5) => fifo_MEMRADDR(5), 
        fifo_MEMRADDR(4) => fifo_MEMRADDR(4), fifo_MEMRADDR(3)
         => fifo_MEMRADDR(3), fifo_MEMRADDR(2) => 
        fifo_MEMRADDR(2), fifo_MEMRADDR(1) => fifo_MEMRADDR(1), 
        fifo_MEMRADDR(0) => fifo_MEMRADDR(0), RDATA_int(7) => 
        RDATA_int(7), RDATA_int(6) => RDATA_int(6), RDATA_int(5)
         => RDATA_int(5), RDATA_int(4) => RDATA_int(4), 
        RDATA_int(3) => RDATA_int(3), RDATA_int(2) => 
        RDATA_int(2), RDATA_int(1) => RDATA_int(1), RDATA_int(0)
         => RDATA_int(0), fifo_MEMWE => fifo_MEMWE, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        fifo_MEMRE => fifo_MEMRE, BIT_CLK => BIT_CLK);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0 is

    port( wptr_bin_sync  : inout std_logic_vector(11 downto 0) := (others => 'Z');
          wptr_gray_sync : in    std_logic_vector(10 downto 0)
        );

end FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0;

architecture DEF_ARCH of 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0 is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    \bin_out_xhdl1_0_a2[1]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(2), B => wptr_bin_sync(3), C
         => wptr_gray_sync(1), Y => wptr_bin_sync(1));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(6), B => wptr_bin_sync(8), C
         => wptr_gray_sync(5), D => wptr_gray_sync(7), Y => 
        wptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(4), B => wptr_gray_sync(3), C
         => wptr_bin_sync(5), D => wptr_gray_sync(2), Y => 
        wptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(2), B => wptr_bin_sync(3), C
         => wptr_gray_sync(0), D => wptr_gray_sync(1), Y => 
        wptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(10), B => wptr_gray_sync(9), Y
         => wptr_bin_sync(9));
    
    \bin_out_xhdl1_i_o2[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(11), B => wptr_gray_sync(10), Y
         => wptr_bin_sync(10));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(7), B => wptr_gray_sync(6), Y
         => wptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(5), B => wptr_gray_sync(4), Y
         => wptr_bin_sync(4));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(9), B => wptr_bin_sync(11), C
         => wptr_gray_sync(8), D => wptr_gray_sync(10), Y => 
        wptr_bin_sync(8));
    
    \bin_out_xhdl1_0_a2[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(8), B => wptr_gray_sync(7), Y
         => wptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(3), B => wptr_gray_sync(4), C
         => wptr_bin_sync(5), Y => wptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1 is

    port( wptr_gray       : in    std_logic_vector(11 downto 0);
          wptr_gray_sync  : out   std_logic_vector(10 downto 0);
          wptr_bin_sync_0 : out   std_logic;
          BIT_CLK         : in    std_logic;
          itx_fifo_rst_i  : in    std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1;

architecture DEF_ARCH of 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \sync_int[10]_net_1\, VCC_net_1, GND_net_1, 
        \sync_int[11]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\, \sync_int[4]_net_1\, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => wptr_gray(9), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => wptr_gray(4), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => wptr_gray(1), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => wptr_gray(11), CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => wptr_gray(6), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_bin_sync_0);
    
    \sync_int[3]\ : SLE
      port map(D => wptr_gray(3), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[3]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => wptr_gray(0), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => wptr_gray(5), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => wptr_gray(2), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => wptr_gray(8), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => wptr_gray(7), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => wptr_gray(10), CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0 is

    port( rptr_gray                 : in    std_logic_vector(11 downto 0);
          rptr_gray_sync            : out   std_logic_vector(10 downto 0);
          rptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          itx_fifo_rst_i            : in    std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0;

architecture DEF_ARCH of 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \sync_int[4]_net_1\, GND_net_1, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\, \sync_int[10]_net_1\, 
        \sync_int[11]_net_1\, \sync_int[1]_net_1\, 
        \sync_int[2]_net_1\, \sync_int[3]_net_1\, 
        \sync_int[0]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => rptr_gray(9), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => rptr_gray(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => rptr_gray(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => rptr_gray(11), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => rptr_gray(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_bin_sync_0);
    
    \sync_int[3]\ : SLE
      port map(D => rptr_gray(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[3]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => rptr_gray(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => rptr_gray(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => rptr_gray(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => rptr_gray(8), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => rptr_gray(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => rptr_gray(10), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv is

    port( rptr_bin_sync  : inout std_logic_vector(11 downto 0) := (others => 'Z');
          rptr_gray_sync : in    std_logic_vector(10 downto 0)
        );

end FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv;

architecture DEF_ARCH of 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    \bin_out_xhdl1_0_a2[1]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(3), B => rptr_gray_sync(1), C
         => rptr_bin_sync(4), D => rptr_gray_sync(2), Y => 
        rptr_bin_sync(1));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(7), B => rptr_gray_sync(6), C
         => rptr_bin_sync(8), D => rptr_gray_sync(5), Y => 
        rptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(4), B => rptr_gray_sync(3), C
         => rptr_gray_sync(2), D => rptr_bin_sync(5), Y => 
        rptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(2), B => rptr_bin_sync(3), C
         => rptr_gray_sync(0), D => rptr_gray_sync(1), Y => 
        rptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2[9]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(10), B => rptr_bin_sync(11), C
         => rptr_gray_sync(9), Y => rptr_bin_sync(9));
    
    \bin_out_xhdl1_i_o2[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(11), B => rptr_gray_sync(10), Y
         => rptr_bin_sync(10));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(8), B => rptr_gray_sync(6), C
         => rptr_gray_sync(7), D => rptr_bin_sync(9), Y => 
        rptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(5), B => rptr_gray_sync(4), C
         => rptr_bin_sync(6), Y => rptr_bin_sync(4));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(10), B => rptr_bin_sync(11), C
         => rptr_gray_sync(9), D => rptr_gray_sync(8), Y => 
        rptr_bin_sync(8));
    
    \bin_out_xhdl1_0_a2[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(8), B => rptr_gray_sync(7), Y
         => rptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(5), B => rptr_gray_sync(4), C
         => rptr_gray_sync(3), D => rptr_bin_sync(6), Y => 
        rptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async is

    port( fifo_MEMWADDR             : out   std_logic_vector(10 downto 0);
          fifo_MEMRADDR             : out   std_logic_vector(10 downto 0);
          TX_FIFO_rd_en             : in    std_logic;
          TX_FIFO_wr_en             : in    std_logic;
          fifo_MEMWE                : out   std_logic;
          fifo_MEMRE                : in    std_logic;
          TX_FIFO_Full              : out   std_logic;
          TX_FIFO_Empty             : out   std_logic;
          un2_re_p                  : in    std_logic;
          BIT_CLK                   : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          itx_fifo_rst_i            : in    std_logic;
          TX_FIFO_OVERFLOW_i        : out   std_logic;
          TX_FIFO_OVERFLOW          : out   std_logic;
          TX_FIFO_UNDERRUN_i        : out   std_logic;
          TX_FIFO_UNDERRUN          : out   std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async;

architecture DEF_ARCH of FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0
    port( wptr_bin_sync  : inout   std_logic_vector(11 downto 0);
          wptr_gray_sync : in    std_logic_vector(10 downto 0) := (others => 'U')
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1
    port( wptr_gray       : in    std_logic_vector(11 downto 0) := (others => 'U');
          wptr_gray_sync  : out   std_logic_vector(10 downto 0);
          wptr_bin_sync_0 : out   std_logic;
          BIT_CLK         : in    std_logic := 'U';
          itx_fifo_rst_i  : in    std_logic := 'U'
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0
    port( rptr_gray                 : in    std_logic_vector(11 downto 0) := (others => 'U');
          rptr_gray_sync            : out   std_logic_vector(10 downto 0);
          rptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          itx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv
    port( rptr_bin_sync  : inout   std_logic_vector(11 downto 0);
          rptr_gray_sync : in    std_logic_vector(10 downto 0) := (others => 'U')
        );
  end component;

    signal \wptr[0]_net_1\, \wptr_s[0]\, \rptr[0]_net_1\, 
        \rptr_s[0]\, \fifo_MEMWADDR[0]\, \memwaddr_r_s[0]\, 
        \fifo_MEMRADDR[0]\, \memraddr_r_s[0]\, \TX_FIFO_UNDERRUN\, 
        \TX_FIFO_OVERFLOW\, \rptr_bin_sync2[10]_net_1\, VCC_net_1, 
        \rptr_bin_sync[10]\, GND_net_1, 
        \rptr_bin_sync2[11]_net_1\, \rptr_bin_sync[11]\, 
        \wptr_gray[0]_net_1\, \wptr_gray_1[0]_net_1\, 
        \wptr_gray[1]_net_1\, \wptr_gray_1[1]_net_1\, 
        \wptr_gray[2]_net_1\, \wptr_gray_1[2]_net_1\, 
        \wptr_gray[3]_net_1\, \wptr_gray_1[3]_net_1\, 
        \wptr_gray[4]_net_1\, \wptr_gray_1[4]_net_1\, 
        \wptr_gray[5]_net_1\, \wptr_gray_1[5]_net_1\, 
        \wptr_gray[6]_net_1\, \wptr_gray_1[6]_net_1\, 
        \wptr_gray[7]_net_1\, \wptr_gray_1[7]_net_1\, 
        \wptr_gray[8]_net_1\, \wptr_gray_1[8]_net_1\, 
        \wptr_gray[9]_net_1\, \wptr_gray_1[9]_net_1\, 
        \wptr_gray[10]_net_1\, \wptr_gray_1[10]_net_1\, 
        \wptr_gray[11]_net_1\, \wptr[11]_net_1\, 
        \wptr_bin_sync2[7]_net_1\, \wptr_bin_sync[7]\, 
        \wptr_bin_sync2[8]_net_1\, \wptr_bin_sync[8]\, 
        \wptr_bin_sync2[9]_net_1\, \wptr_bin_sync[9]\, 
        \wptr_bin_sync2[10]_net_1\, \wptr_bin_sync[10]\, 
        \wptr_bin_sync2[11]_net_1\, \wptr_bin_sync[11]\, 
        \rptr_bin_sync2[0]_net_1\, \rptr_bin_sync[0]\, 
        \rptr_bin_sync2[1]_net_1\, \rptr_bin_sync[1]\, 
        \rptr_bin_sync2[2]_net_1\, \rptr_bin_sync[2]\, 
        \rptr_bin_sync2[3]_net_1\, \rptr_bin_sync[3]\, 
        \rptr_bin_sync2[4]_net_1\, \rptr_bin_sync[4]\, 
        \rptr_bin_sync2[5]_net_1\, \rptr_bin_sync[5]\, 
        \rptr_bin_sync2[6]_net_1\, \rptr_bin_sync[6]\, 
        \rptr_bin_sync2[7]_net_1\, \rptr_bin_sync[7]\, 
        \rptr_bin_sync2[8]_net_1\, \rptr_bin_sync[8]\, 
        \rptr_bin_sync2[9]_net_1\, \rptr_bin_sync[9]\, rdiff_bus, 
        \wptr_bin_sync[0]\, \wptr_bin_sync2[1]_net_1\, 
        \wptr_bin_sync[1]\, \wptr_bin_sync2[2]_net_1\, 
        \wptr_bin_sync[2]\, \wptr_bin_sync2[3]_net_1\, 
        \wptr_bin_sync[3]\, \wptr_bin_sync2[4]_net_1\, 
        \wptr_bin_sync[4]\, \wptr_bin_sync2[5]_net_1\, 
        \wptr_bin_sync[5]\, \wptr_bin_sync2[6]_net_1\, 
        \wptr_bin_sync[6]\, \rptr_gray[7]_net_1\, 
        \rptr_gray_1[7]_net_1\, \rptr_gray[8]_net_1\, 
        \rptr_gray_1[8]_net_1\, \rptr_gray[9]_net_1\, 
        \rptr_gray_1[9]_net_1\, \rptr_gray[10]_net_1\, 
        \rptr_gray_1[10]_net_1\, \rptr_gray[11]_net_1\, 
        \rptr[11]_net_1\, \rptr_gray[0]_net_1\, 
        \rptr_gray_1[0]_net_1\, \rptr_gray[1]_net_1\, 
        \rptr_gray_1[1]_net_1\, \rptr_gray[2]_net_1\, 
        \rptr_gray_1[2]_net_1\, \rptr_gray[3]_net_1\, 
        \rptr_gray_1[3]_net_1\, \rptr_gray[4]_net_1\, 
        \rptr_gray_1[4]_net_1\, \rptr_gray[5]_net_1\, 
        \rptr_gray_1[5]_net_1\, \rptr_gray[6]_net_1\, 
        \rptr_gray_1[6]_net_1\, un1_we_p, empty_r_3, 
        \TX_FIFO_Full\, \fulli\, \fifo_MEMRADDR[1]\, 
        \memraddr_r_s[1]\, \fifo_MEMRADDR[2]\, \memraddr_r_s[2]\, 
        \fifo_MEMRADDR[3]\, \memraddr_r_s[3]\, \fifo_MEMRADDR[4]\, 
        \memraddr_r_s[4]\, \fifo_MEMRADDR[5]\, \memraddr_r_s[5]\, 
        \fifo_MEMRADDR[6]\, \memraddr_r_s[6]\, \fifo_MEMRADDR[7]\, 
        \memraddr_r_s[7]\, \fifo_MEMRADDR[8]\, \memraddr_r_s[8]\, 
        \fifo_MEMRADDR[9]\, \memraddr_r_s[9]\, 
        \fifo_MEMRADDR[10]\, \memraddr_r_s[10]_net_1\, 
        \fifo_MEMWE\, \fifo_MEMWADDR[1]\, \memwaddr_r_s[1]\, 
        \fifo_MEMWADDR[2]\, \memwaddr_r_s[2]\, \fifo_MEMWADDR[3]\, 
        \memwaddr_r_s[3]\, \fifo_MEMWADDR[4]\, \memwaddr_r_s[4]\, 
        \fifo_MEMWADDR[5]\, \memwaddr_r_s[5]\, \fifo_MEMWADDR[6]\, 
        \memwaddr_r_s[6]\, \fifo_MEMWADDR[7]\, \memwaddr_r_s[7]\, 
        \fifo_MEMWADDR[8]\, \memwaddr_r_s[8]\, \fifo_MEMWADDR[9]\, 
        \memwaddr_r_s[9]\, \fifo_MEMWADDR[10]\, 
        \memwaddr_r_s[10]_net_1\, \rptr[1]_net_1\, \rptr_s[1]\, 
        \rptr[2]_net_1\, \rptr_s[2]\, \rptr[3]_net_1\, 
        \rptr_s[3]\, \rptr[4]_net_1\, \rptr_s[4]\, 
        \rptr[5]_net_1\, \rptr_s[5]\, \rptr[6]_net_1\, 
        \rptr_s[6]\, \rptr[7]_net_1\, \rptr_s[7]\, 
        \rptr[8]_net_1\, \rptr_s[8]\, \rptr[9]_net_1\, 
        \rptr_s[9]\, \rptr[10]_net_1\, \rptr_s[10]\, 
        \rptr_s[11]_net_1\, \wptr[1]_net_1\, \wptr_s[1]\, 
        \wptr[2]_net_1\, \wptr_s[2]\, \wptr[3]_net_1\, 
        \wptr_s[3]\, \wptr[4]_net_1\, \wptr_s[4]\, 
        \wptr[5]_net_1\, \wptr_s[5]\, \wptr[6]_net_1\, 
        \wptr_s[6]\, \wptr[7]_net_1\, \wptr_s[7]\, 
        \wptr[8]_net_1\, \wptr_s[8]\, \wptr[9]_net_1\, 
        \wptr_s[9]\, \wptr[10]_net_1\, \wptr_s[10]\, 
        \wptr_s[11]_net_1\, \wdiff_bus_cry_0\, wdiff_bus_cry_0_Y, 
        \wdiff_bus_cry_1\, \wdiff_bus[1]\, \wdiff_bus_cry_2\, 
        \wdiff_bus[2]\, \wdiff_bus_cry_3\, \wdiff_bus[3]\, 
        \wdiff_bus_cry_4\, \wdiff_bus[4]\, \wdiff_bus_cry_5\, 
        \wdiff_bus[5]\, \wdiff_bus_cry_6\, \wdiff_bus[6]\, 
        \wdiff_bus_cry_7\, \wdiff_bus[7]\, \wdiff_bus_cry_8\, 
        \wdiff_bus[8]\, \wdiff_bus_cry_9\, \wdiff_bus[9]\, 
        \wdiff_bus[11]\, \wdiff_bus_cry_10\, \wdiff_bus[10]\, 
        \rdiff_bus_cry_0\, rdiff_bus_cry_0_Y, \rdiff_bus_cry_1\, 
        \rdiff_bus[1]\, \rdiff_bus_cry_2\, \rdiff_bus[2]\, 
        \rdiff_bus_cry_3\, \rdiff_bus[3]\, \rdiff_bus_cry_4\, 
        \rdiff_bus[4]\, \rdiff_bus_cry_5\, \rdiff_bus[5]\, 
        \rdiff_bus_cry_6\, \rdiff_bus[6]\, \rdiff_bus_cry_7\, 
        \rdiff_bus[7]\, \rdiff_bus_cry_8\, \rdiff_bus[8]\, 
        \rdiff_bus_cry_9\, \rdiff_bus[9]\, \rdiff_bus[11]\, 
        \rdiff_bus_cry_10\, \rdiff_bus[10]\, wptr_s_267_FCO, 
        \wptr_cry[1]_net_1\, \wptr_cry[2]_net_1\, 
        \wptr_cry[3]_net_1\, \wptr_cry[4]_net_1\, 
        \wptr_cry[5]_net_1\, \wptr_cry[6]_net_1\, 
        \wptr_cry[7]_net_1\, \wptr_cry[8]_net_1\, 
        \wptr_cry[9]_net_1\, \wptr_cry[10]_net_1\, rptr_s_268_FCO, 
        \rptr_cry[1]_net_1\, \rptr_cry[2]_net_1\, 
        \rptr_cry[3]_net_1\, \rptr_cry[4]_net_1\, 
        \rptr_cry[5]_net_1\, \rptr_cry[6]_net_1\, 
        \rptr_cry[7]_net_1\, \rptr_cry[8]_net_1\, 
        \rptr_cry[9]_net_1\, \rptr_cry[10]_net_1\, 
        memwaddr_r_s_269_FCO, \memwaddr_r_cry[1]_net_1\, 
        \memwaddr_r_cry[2]_net_1\, \memwaddr_r_cry[3]_net_1\, 
        \memwaddr_r_cry[4]_net_1\, \memwaddr_r_cry[5]_net_1\, 
        \memwaddr_r_cry[6]_net_1\, \memwaddr_r_cry[7]_net_1\, 
        \memwaddr_r_cry[8]_net_1\, \memwaddr_r_cry[9]_net_1\, 
        memraddr_r_s_270_FCO, \memraddr_r_cry[1]_net_1\, 
        \memraddr_r_cry[2]_net_1\, \memraddr_r_cry[3]_net_1\, 
        \memraddr_r_cry[4]_net_1\, \memraddr_r_cry[5]_net_1\, 
        \memraddr_r_cry[6]_net_1\, \memraddr_r_cry[7]_net_1\, 
        \memraddr_r_cry[8]_net_1\, \memraddr_r_cry[9]_net_1\, 
        empty_r_3_0_a2_1, empty_r_3_0_a2_7, un4_fullilto10_i_a2_7, 
        un4_fullilto10_i_a2_6, empty_r_3_0_a2_9, empty_r_3_0_a2_5, 
        un4_fullilto10_i_a2_8, \wptr_gray_sync[0]\, 
        \wptr_gray_sync[1]\, \wptr_gray_sync[2]\, 
        \wptr_gray_sync[3]\, \wptr_gray_sync[4]\, 
        \wptr_gray_sync[5]\, \wptr_gray_sync[6]\, 
        \wptr_gray_sync[7]\, \wptr_gray_sync[8]\, 
        \wptr_gray_sync[9]\, \wptr_gray_sync[10]\, 
        \rptr_gray_sync[0]\, \rptr_gray_sync[1]\, 
        \rptr_gray_sync[2]\, \rptr_gray_sync[3]\, 
        \rptr_gray_sync[4]\, \rptr_gray_sync[5]\, 
        \rptr_gray_sync[6]\, \rptr_gray_sync[7]\, 
        \rptr_gray_sync[8]\, \rptr_gray_sync[9]\, 
        \rptr_gray_sync[10]\ : std_logic;

    for all : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0
	Use entity work.
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0(DEF_ARCH);
    for all : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1
	Use entity work.
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1(DEF_ARCH);
    for all : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0
	Use entity work.
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0(DEF_ARCH);
    for all : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv
	Use entity work.
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv(DEF_ARCH);
begin 

    fifo_MEMWADDR(10) <= \fifo_MEMWADDR[10]\;
    fifo_MEMWADDR(9) <= \fifo_MEMWADDR[9]\;
    fifo_MEMWADDR(8) <= \fifo_MEMWADDR[8]\;
    fifo_MEMWADDR(7) <= \fifo_MEMWADDR[7]\;
    fifo_MEMWADDR(6) <= \fifo_MEMWADDR[6]\;
    fifo_MEMWADDR(5) <= \fifo_MEMWADDR[5]\;
    fifo_MEMWADDR(4) <= \fifo_MEMWADDR[4]\;
    fifo_MEMWADDR(3) <= \fifo_MEMWADDR[3]\;
    fifo_MEMWADDR(2) <= \fifo_MEMWADDR[2]\;
    fifo_MEMWADDR(1) <= \fifo_MEMWADDR[1]\;
    fifo_MEMWADDR(0) <= \fifo_MEMWADDR[0]\;
    fifo_MEMRADDR(10) <= \fifo_MEMRADDR[10]\;
    fifo_MEMRADDR(9) <= \fifo_MEMRADDR[9]\;
    fifo_MEMRADDR(8) <= \fifo_MEMRADDR[8]\;
    fifo_MEMRADDR(7) <= \fifo_MEMRADDR[7]\;
    fifo_MEMRADDR(6) <= \fifo_MEMRADDR[6]\;
    fifo_MEMRADDR(5) <= \fifo_MEMRADDR[5]\;
    fifo_MEMRADDR(4) <= \fifo_MEMRADDR[4]\;
    fifo_MEMRADDR(3) <= \fifo_MEMRADDR[3]\;
    fifo_MEMRADDR(2) <= \fifo_MEMRADDR[2]\;
    fifo_MEMRADDR(1) <= \fifo_MEMRADDR[1]\;
    fifo_MEMRADDR(0) <= \fifo_MEMRADDR[0]\;
    fifo_MEMWE <= \fifo_MEMWE\;
    TX_FIFO_Full <= \TX_FIFO_Full\;
    TX_FIFO_OVERFLOW <= \TX_FIFO_OVERFLOW\;
    TX_FIFO_UNDERRUN <= \TX_FIFO_UNDERRUN\;

    \rptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[4]_net_1\, S
         => \rptr_s[5]\, Y => OPEN, FCO => \rptr_cry[5]_net_1\);
    
    underflow_r_RNIFFTA : CFG1
      generic map(INIT => "01")

      port map(A => \TX_FIFO_UNDERRUN\, Y => TX_FIFO_UNDERRUN_i);
    
    wdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[8]_net_1\, B => 
        \rptr_bin_sync2[8]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_7\, S => \wdiff_bus[8]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_8\);
    
    \wptr_gray[4]\ : SLE
      port map(D => \wptr_gray_1[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[4]_net_1\);
    
    \rptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[3]_net_1\, B => \rptr[4]_net_1\, Y => 
        \rptr_gray_1[3]_net_1\);
    
    \rptr_bin_sync2[6]\ : SLE
      port map(D => \rptr_bin_sync[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[6]_net_1\);
    
    \rptr[1]\ : SLE
      port map(D => \rptr_s[1]\, CLK => BIT_CLK, EN => fifo_MEMRE, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[1]_net_1\);
    
    \wptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[9]_net_1\, B => \wptr[10]_net_1\, Y => 
        \wptr_gray_1[9]_net_1\);
    
    \rptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[5]_net_1\, B => \rptr[6]_net_1\, Y => 
        \rptr_gray_1[5]_net_1\);
    
    \rptr_gray[9]\ : SLE
      port map(D => \rptr_gray_1[9]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[9]_net_1\);
    
    \rptr_gray[8]\ : SLE
      port map(D => \rptr_gray_1[8]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[8]_net_1\);
    
    \rptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[2]_net_1\, B => \rptr[3]_net_1\, Y => 
        \rptr_gray_1[2]_net_1\);
    
    \rptr_bin_sync2[7]\ : SLE
      port map(D => \rptr_bin_sync[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[7]_net_1\);
    
    \memwaddr_r[1]\ : SLE
      port map(D => \memwaddr_r_s[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[1]\);
    
    fulli : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \wdiff_bus[11]\, B => TX_FIFO_wr_en, C => 
        un4_fullilto10_i_a2_8, D => un4_fullilto10_i_a2_7, Y => 
        \fulli\);
    
    \memwaddr_r_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[5]_net_1\, S => \memwaddr_r_s[6]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[6]_net_1\);
    
    \memwaddr_r_s[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[9]_net_1\, S => \memwaddr_r_s[10]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \wptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[7]_net_1\, B => \wptr[8]_net_1\, Y => 
        \wptr_gray_1[7]_net_1\);
    
    \memraddr_r[0]\ : SLE
      port map(D => \memraddr_r_s[0]\, CLK => BIT_CLK, EN => 
        fifo_MEMRE, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[0]\);
    
    \wptr[0]\ : SLE
      port map(D => \wptr_s[0]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[0]_net_1\);
    
    \rptr_bin_sync2[8]\ : SLE
      port map(D => \rptr_bin_sync[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[8]_net_1\);
    
    \rptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[1]_net_1\, B => \rptr[2]_net_1\, Y => 
        \rptr_gray_1[1]_net_1\);
    
    \rptr_gray[10]\ : SLE
      port map(D => \rptr_gray_1[10]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[10]_net_1\);
    
    \wptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[0]_net_1\, B => \wptr[1]_net_1\, Y => 
        \wptr_gray_1[0]_net_1\);
    
    wdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[9]_net_1\, B => 
        \rptr_bin_sync2[9]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_8\, S => \wdiff_bus[9]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_9\);
    
    \rptr[5]\ : SLE
      port map(D => \rptr_s[5]\, CLK => BIT_CLK, EN => fifo_MEMRE, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[5]_net_1\);
    
    \rptr_gray[3]\ : SLE
      port map(D => \rptr_gray_1[3]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[3]_net_1\);
    
    \rptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[5]_net_1\, S
         => \rptr_s[6]\, Y => OPEN, FCO => \rptr_cry[6]_net_1\);
    
    \memwaddr_r_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => memwaddr_r_s_269_FCO, S
         => \memwaddr_r_s[1]\, Y => OPEN, FCO => 
        \memwaddr_r_cry[1]_net_1\);
    
    \wptr_gray[3]\ : SLE
      port map(D => \wptr_gray_1[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[3]_net_1\);
    
    \rptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[11]_net_1\, B => \rptr[10]_net_1\, Y
         => \rptr_gray_1[10]_net_1\);
    
    wdiff_bus_s_11 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr_bin_sync2[11]_net_1\, C
         => \wptr[11]_net_1\, D => GND_net_1, FCI => 
        \wdiff_bus_cry_10\, S => \wdiff_bus[11]\, Y => OPEN, FCO
         => OPEN);
    
    \rptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[7]_net_1\, S
         => \rptr_s[8]\, Y => OPEN, FCO => \rptr_cry[8]_net_1\);
    
    \rptr[7]\ : SLE
      port map(D => \rptr_s[7]\, CLK => BIT_CLK, EN => fifo_MEMRE, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[7]_net_1\);
    
    rdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[4]_net_1\, B => 
        \rptr[4]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_3\, S => \rdiff_bus[4]\, Y => OPEN, FCO
         => \rdiff_bus_cry_4\);
    
    \rptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[9]_net_1\, S
         => \rptr_s[10]\, Y => OPEN, FCO => \rptr_cry[10]_net_1\);
    
    \rptr_bin_sync2[0]\ : SLE
      port map(D => \rptr_bin_sync[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[0]_net_1\);
    
    \L1.empty_r_3_0_a2_7\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \rdiff_bus[5]\, B => \rdiff_bus[6]\, C => 
        \rdiff_bus[7]\, D => \rdiff_bus[8]\, Y => 
        empty_r_3_0_a2_7);
    
    \wptr[11]\ : SLE
      port map(D => \wptr_s[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \wptr[11]_net_1\);
    
    rdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[1]_net_1\, B => 
        \rptr[1]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_0\, S => \rdiff_bus[1]\, Y => OPEN, FCO
         => \rdiff_bus_cry_1\);
    
    \memraddr_r[1]\ : SLE
      port map(D => \memraddr_r_s[1]\, CLK => BIT_CLK, EN => 
        fifo_MEMRE, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[1]\);
    
    \L1.empty_r_3_0_a2_9\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \rdiff_bus[1]\, B => \rdiff_bus[2]\, C => 
        empty_r_3_0_a2_7, D => empty_r_3_0_a2_1, Y => 
        empty_r_3_0_a2_9);
    
    rptr_s_268 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => rptr_s_268_FCO);
    
    \rptr_bin_sync2[2]\ : SLE
      port map(D => \rptr_bin_sync[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[2]_net_1\);
    
    rdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[6]_net_1\, B => 
        \rptr[6]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_5\, S => \rdiff_bus[6]\, Y => OPEN, FCO
         => \rdiff_bus_cry_6\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \memwaddr_r_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[2]_net_1\, S => \memwaddr_r_s[3]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[3]_net_1\);
    
    \rptr_gray[1]\ : SLE
      port map(D => \rptr_gray_1[1]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[1]_net_1\);
    
    \memwaddr_r[7]\ : SLE
      port map(D => \memwaddr_r_s[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[7]\);
    
    \memraddr_r_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[1]_net_1\, S => \memraddr_r_s[2]\, Y => 
        OPEN, FCO => \memraddr_r_cry[2]_net_1\);
    
    \wptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[3]_net_1\, S
         => \wptr_s[4]\, Y => OPEN, FCO => \wptr_cry[4]_net_1\);
    
    \memraddr_r_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[7]_net_1\, S => \memraddr_r_s[8]\, Y => 
        OPEN, FCO => \memraddr_r_cry[8]_net_1\);
    
    \wptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[9]_net_1\, S
         => \wptr_s[10]\, Y => OPEN, FCO => \wptr_cry[10]_net_1\);
    
    wdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[5]_net_1\, B => 
        \rptr_bin_sync2[5]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_4\, S => \wdiff_bus[5]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_5\);
    
    \memwaddr_r[4]\ : SLE
      port map(D => \memwaddr_r_s[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[4]\);
    
    \wptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[1]_net_1\, S
         => \wptr_s[2]\, Y => OPEN, FCO => \wptr_cry[2]_net_1\);
    
    wdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[0]_net_1\, B => 
        \rptr_bin_sync2[0]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => VCC_net_1, S => OPEN, Y => wdiff_bus_cry_0_Y, FCO
         => \wdiff_bus_cry_0\);
    
    \wptr[1]\ : SLE
      port map(D => \wptr_s[1]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[1]_net_1\);
    
    \rptr_bin_sync2[4]\ : SLE
      port map(D => \rptr_bin_sync[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[4]_net_1\);
    
    \wptr_bin_sync2[6]\ : SLE
      port map(D => \wptr_bin_sync[6]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[6]_net_1\);
    
    \L1.un1_we_p\ : CFG2
      generic map(INIT => x"8")

      port map(A => \TX_FIFO_Full\, B => TX_FIFO_wr_en, Y => 
        un1_we_p);
    
    \rptr[3]\ : SLE
      port map(D => \rptr_s[3]\, CLK => BIT_CLK, EN => fifo_MEMRE, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[3]_net_1\);
    
    \wptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[2]_net_1\, S
         => \wptr_s[3]\, Y => OPEN, FCO => \wptr_cry[3]_net_1\);
    
    \rptr[6]\ : SLE
      port map(D => \rptr_s[6]\, CLK => BIT_CLK, EN => fifo_MEMRE, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[6]_net_1\);
    
    rdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[8]_net_1\, B => 
        \rptr[8]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_7\, S => \rdiff_bus[8]\, Y => OPEN, FCO
         => \rdiff_bus_cry_8\);
    
    \wptr_gray[10]\ : SLE
      port map(D => \wptr_gray_1[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[10]_net_1\);
    
    rdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[7]_net_1\, B => 
        \rptr[7]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_6\, S => \rdiff_bus[7]\, Y => OPEN, FCO
         => \rdiff_bus_cry_7\);
    
    \wptr_bin_sync2[7]\ : SLE
      port map(D => \wptr_bin_sync[7]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[7]_net_1\);
    
    overflow_r_RNIDBD3 : CFG1
      generic map(INIT => "01")

      port map(A => \TX_FIFO_OVERFLOW\, Y => TX_FIFO_OVERFLOW_i);
    
    \rptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[8]_net_1\, S
         => \rptr_s[9]\, Y => OPEN, FCO => \rptr_cry[9]_net_1\);
    
    \T11.un4_fullilto10_i_a2_8\ : CFG4
      generic map(INIT => x"4000")

      port map(A => wdiff_bus_cry_0_Y, B => \wdiff_bus[1]\, C => 
        \wdiff_bus[10]\, D => un4_fullilto10_i_a2_6, Y => 
        un4_fullilto10_i_a2_8);
    
    \rptr_gray[5]\ : SLE
      port map(D => \rptr_gray_1[5]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[5]_net_1\);
    
    \wptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[2]_net_1\, B => \wptr[3]_net_1\, Y => 
        \wptr_gray_1[2]_net_1\);
    
    \wptr[5]\ : SLE
      port map(D => \wptr_s[5]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[5]_net_1\);
    
    rdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[5]_net_1\, B => 
        \rptr[5]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_4\, S => \rdiff_bus[5]\, Y => OPEN, FCO
         => \rdiff_bus_cry_5\);
    
    \wptr_bin_sync2[8]\ : SLE
      port map(D => \wptr_bin_sync[8]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[8]_net_1\);
    
    \wptr[7]\ : SLE
      port map(D => \wptr_s[7]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[7]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \wptr_gray[1]\ : SLE
      port map(D => \wptr_gray_1[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[1]_net_1\);
    
    \rptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[9]_net_1\, B => \rptr[10]_net_1\, Y => 
        \rptr_gray_1[9]_net_1\);
    
    \rptr_bin_sync2[5]\ : SLE
      port map(D => \rptr_bin_sync[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[5]_net_1\);
    
    \rptr_bin_sync2[1]\ : SLE
      port map(D => \rptr_bin_sync[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[1]_net_1\);
    
    \memwaddr_r[10]\ : SLE
      port map(D => \memwaddr_r_s[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[10]\);
    
    wdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[7]_net_1\, B => 
        \rptr_bin_sync2[7]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_6\, S => \wdiff_bus[7]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_7\);
    
    \wptr_bin_sync2[0]\ : SLE
      port map(D => \wptr_bin_sync[0]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        rdiff_bus);
    
    \L1.empty_r_3_0_a2_1\ : CFG2
      generic map(INIT => x"1")

      port map(A => \rdiff_bus[4]\, B => \rdiff_bus[3]\, Y => 
        empty_r_3_0_a2_1);
    
    rdiff_bus_s_11 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        \wptr_bin_sync2[11]_net_1\, D => GND_net_1, FCI => 
        \rdiff_bus_cry_10\, S => \rdiff_bus[11]\, Y => OPEN, FCO
         => OPEN);
    
    \memwaddr_r_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[7]_net_1\, S => \memwaddr_r_s[8]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[8]_net_1\);
    
    \wptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => wptr_s_267_FCO, S => 
        \wptr_s[1]\, Y => OPEN, FCO => \wptr_cry[1]_net_1\);
    
    \memraddr_r[8]\ : SLE
      port map(D => \memraddr_r_s[8]\, CLK => BIT_CLK, EN => 
        fifo_MEMRE, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[8]\);
    
    \rptr[9]\ : SLE
      port map(D => \rptr_s[9]\, CLK => BIT_CLK, EN => fifo_MEMRE, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[9]_net_1\);
    
    \wptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[6]_net_1\, B => \wptr[7]_net_1\, Y => 
        \wptr_gray_1[6]_net_1\);
    
    \wptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[6]_net_1\, S
         => \wptr_s[7]\, Y => OPEN, FCO => \wptr_cry[7]_net_1\);
    
    \wptr_bin_sync2[2]\ : SLE
      port map(D => \wptr_bin_sync[2]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[2]_net_1\);
    
    \T11.un4_fullilto10_i_a2_6\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[2]\, B => \wdiff_bus[3]\, C => 
        \wdiff_bus[5]\, D => \wdiff_bus[4]\, Y => 
        un4_fullilto10_i_a2_6);
    
    \rptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \rptr[0]_net_1\, Y => \rptr_s[0]\);
    
    \rptr[4]\ : SLE
      port map(D => \rptr_s[4]\, CLK => BIT_CLK, EN => fifo_MEMRE, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[4]_net_1\);
    
    \memwaddr_r_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[4]_net_1\, S => \memwaddr_r_s[5]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[5]_net_1\);
    
    \memraddr_r_s[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[9]_net_1\, S => \memraddr_r_s[10]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \wptr_gray[6]\ : SLE
      port map(D => \wptr_gray_1[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[6]_net_1\);
    
    \wptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[3]_net_1\, B => \wptr[4]_net_1\, Y => 
        \wptr_gray_1[3]_net_1\);
    
    \wptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[4]_net_1\, S
         => \wptr_s[5]\, Y => OPEN, FCO => \wptr_cry[5]_net_1\);
    
    \memraddr_r_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[4]_net_1\, S => \memraddr_r_s[5]\, Y => 
        OPEN, FCO => \memraddr_r_cry[5]_net_1\);
    
    \memraddr_r_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => memraddr_r_s_270_FCO, S
         => \memraddr_r_s[1]\, Y => OPEN, FCO => 
        \memraddr_r_cry[1]_net_1\);
    
    \rptr_gray[4]\ : SLE
      port map(D => \rptr_gray_1[4]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[4]_net_1\);
    
    \wptr_bin_sync2[4]\ : SLE
      port map(D => \wptr_bin_sync[4]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[4]_net_1\);
    
    \wptr[3]\ : SLE
      port map(D => \wptr_s[3]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[3]_net_1\);
    
    \memwaddr_r[6]\ : SLE
      port map(D => \memwaddr_r_s[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[6]\);
    
    \wptr_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[10]_net_1\, S
         => \wptr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \wptr[6]\ : SLE
      port map(D => \wptr_s[6]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[6]_net_1\);
    
    \memwaddr_r[9]\ : SLE
      port map(D => \memwaddr_r_s[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[9]\);
    
    \memraddr_r_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[3]_net_1\, S => \memraddr_r_s[4]\, Y => 
        OPEN, FCO => \memraddr_r_cry[4]_net_1\);
    
    \memraddr_r[10]\ : SLE
      port map(D => \memraddr_r_s[10]_net_1\, CLK => BIT_CLK, EN
         => fifo_MEMRE, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \fifo_MEMRADDR[10]\);
    
    \memwaddr_r[3]\ : SLE
      port map(D => \memwaddr_r_s[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[3]\);
    
    full_r : SLE
      port map(D => \fulli\, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \TX_FIFO_Full\);
    
    \rptr_bin_sync2[3]\ : SLE
      port map(D => \rptr_bin_sync[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[3]_net_1\);
    
    \wptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \wptr[0]_net_1\, Y => \wptr_s[0]\);
    
    \rptr[2]\ : SLE
      port map(D => \rptr_s[2]\, CLK => BIT_CLK, EN => fifo_MEMRE, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[2]_net_1\);
    
    \memraddr_r[3]\ : SLE
      port map(D => \memraddr_r_s[3]\, CLK => BIT_CLK, EN => 
        fifo_MEMRE, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[3]\);
    
    \rptr_bin_sync2[9]\ : SLE
      port map(D => \rptr_bin_sync[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[9]_net_1\);
    
    \rptr[11]\ : SLE
      port map(D => \rptr_s[11]_net_1\, CLK => BIT_CLK, EN => 
        fifo_MEMRE, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rptr[11]_net_1\);
    
    \wptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[5]_net_1\, S
         => \wptr_s[6]\, Y => OPEN, FCO => \wptr_cry[6]_net_1\);
    
    \rptr_bin_sync2[11]\ : SLE
      port map(D => \rptr_bin_sync[11]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[11]_net_1\);
    
    \wptr_bin_sync2[5]\ : SLE
      port map(D => \wptr_bin_sync[5]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[5]_net_1\);
    
    \wptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[7]_net_1\, S
         => \wptr_s[8]\, Y => OPEN, FCO => \wptr_cry[8]_net_1\);
    
    \wptr_bin_sync2[1]\ : SLE
      port map(D => \wptr_bin_sync[1]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[1]_net_1\);
    
    Wr_corefifo_grayToBinConv : 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0
      port map(wptr_bin_sync(11) => \wptr_bin_sync[11]\, 
        wptr_bin_sync(10) => \wptr_bin_sync[10]\, 
        wptr_bin_sync(9) => \wptr_bin_sync[9]\, wptr_bin_sync(8)
         => \wptr_bin_sync[8]\, wptr_bin_sync(7) => 
        \wptr_bin_sync[7]\, wptr_bin_sync(6) => 
        \wptr_bin_sync[6]\, wptr_bin_sync(5) => 
        \wptr_bin_sync[5]\, wptr_bin_sync(4) => 
        \wptr_bin_sync[4]\, wptr_bin_sync(3) => 
        \wptr_bin_sync[3]\, wptr_bin_sync(2) => 
        \wptr_bin_sync[2]\, wptr_bin_sync(1) => 
        \wptr_bin_sync[1]\, wptr_bin_sync(0) => 
        \wptr_bin_sync[0]\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\);
    
    \wptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[4]_net_1\, B => \wptr[5]_net_1\, Y => 
        \wptr_gray_1[4]_net_1\);
    
    overflow_r : SLE
      port map(D => un1_we_p, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \TX_FIFO_OVERFLOW\);
    
    \memraddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMRADDR[0]\, Y => \memraddr_r_s[0]\);
    
    \rptr_gray[11]\ : SLE
      port map(D => \rptr[11]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[10]\ : SLE
      port map(D => \wptr_bin_sync[10]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[10]_net_1\);
    
    \rptr[10]\ : SLE
      port map(D => \rptr_s[10]\, CLK => BIT_CLK, EN => 
        fifo_MEMRE, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rptr[10]_net_1\);
    
    \wptr[9]\ : SLE
      port map(D => \wptr_s[9]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[9]_net_1\);
    
    Wr_corefifo_doubleSync : 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1
      port map(wptr_gray(11) => \wptr_gray[11]_net_1\, 
        wptr_gray(10) => \wptr_gray[10]_net_1\, wptr_gray(9) => 
        \wptr_gray[9]_net_1\, wptr_gray(8) => 
        \wptr_gray[8]_net_1\, wptr_gray(7) => 
        \wptr_gray[7]_net_1\, wptr_gray(6) => 
        \wptr_gray[6]_net_1\, wptr_gray(5) => 
        \wptr_gray[5]_net_1\, wptr_gray(4) => 
        \wptr_gray[4]_net_1\, wptr_gray(3) => 
        \wptr_gray[3]_net_1\, wptr_gray(2) => 
        \wptr_gray[2]_net_1\, wptr_gray(1) => 
        \wptr_gray[1]_net_1\, wptr_gray(0) => 
        \wptr_gray[0]_net_1\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\, wptr_bin_sync_0 => 
        \wptr_bin_sync[11]\, BIT_CLK => BIT_CLK, itx_fifo_rst_i
         => itx_fifo_rst_i);
    
    \rptr_gray[0]\ : SLE
      port map(D => \rptr_gray_1[0]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[0]_net_1\);
    
    empty_r : SLE
      port map(D => empty_r_3, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => TX_FIFO_Empty);
    
    \memwaddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMWADDR[0]\, Y => \memwaddr_r_s[0]\);
    
    \T11.un4_fullilto10_i_a2_7\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[6]\, B => \wdiff_bus[7]\, C => 
        \wdiff_bus[8]\, D => \wdiff_bus[9]\, Y => 
        un4_fullilto10_i_a2_7);
    
    \rptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[7]_net_1\, B => \rptr[8]_net_1\, Y => 
        \rptr_gray_1[7]_net_1\);
    
    \wptr[4]\ : SLE
      port map(D => \wptr_s[4]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[4]_net_1\);
    
    \memwaddr_r[8]\ : SLE
      port map(D => \memwaddr_r_s[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[8]\);
    
    \memwaddr_r[2]\ : SLE
      port map(D => \memwaddr_r_s[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[2]\);
    
    \L1.empty_r_3_0_a2_5\ : CFG3
      generic map(INIT => x"54")

      port map(A => \rdiff_bus[11]\, B => TX_FIFO_rd_en, C => 
        rdiff_bus_cry_0_Y, Y => empty_r_3_0_a2_5);
    
    \wptr_bin_sync2[11]\ : SLE
      port map(D => \wptr_bin_sync[11]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[11]_net_1\);
    
    memwe : CFG2
      generic map(INIT => x"4")

      port map(A => \TX_FIFO_Full\, B => TX_FIFO_wr_en, Y => 
        \fifo_MEMWE\);
    
    \wptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[1]_net_1\, B => \wptr[2]_net_1\, Y => 
        \wptr_gray_1[1]_net_1\);
    
    underflow_r : SLE
      port map(D => un2_re_p, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_UNDERRUN\);
    
    \memwaddr_r_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[6]_net_1\, S => \memwaddr_r_s[7]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[7]_net_1\);
    
    \wptr_gray[5]\ : SLE
      port map(D => \wptr_gray_1[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[5]_net_1\);
    
    \memraddr_r[7]\ : SLE
      port map(D => \memraddr_r_s[7]\, CLK => BIT_CLK, EN => 
        fifo_MEMRE, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[7]\);
    
    \rptr_bin_sync2[10]\ : SLE
      port map(D => \rptr_bin_sync[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[10]_net_1\);
    
    wdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[10]_net_1\, B => 
        \rptr_bin_sync2[10]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_9\, S => \wdiff_bus[10]\, 
        Y => OPEN, FCO => \wdiff_bus_cry_10\);
    
    \memwaddr_r_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[8]_net_1\, S => \memwaddr_r_s[9]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[9]_net_1\);
    
    \wptr_gray[8]\ : SLE
      port map(D => \wptr_gray_1[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[8]_net_1\);
    
    \wptr_gray[7]\ : SLE
      port map(D => \wptr_gray_1[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[7]_net_1\);
    
    \wptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[5]_net_1\, B => \wptr[6]_net_1\, Y => 
        \wptr_gray_1[5]_net_1\);
    
    \memwaddr_r[5]\ : SLE
      port map(D => \memwaddr_r_s[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[5]\);
    
    \L1.empty_r_3_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \rdiff_bus[9]\, B => \rdiff_bus[10]\, C => 
        empty_r_3_0_a2_5, D => empty_r_3_0_a2_9, Y => empty_r_3);
    
    \rptr[8]\ : SLE
      port map(D => \rptr_s[8]\, CLK => BIT_CLK, EN => fifo_MEMRE, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[8]_net_1\);
    
    Rd_corefifo_doubleSync : 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0
      port map(rptr_gray(11) => \rptr_gray[11]_net_1\, 
        rptr_gray(10) => \rptr_gray[10]_net_1\, rptr_gray(9) => 
        \rptr_gray[9]_net_1\, rptr_gray(8) => 
        \rptr_gray[8]_net_1\, rptr_gray(7) => 
        \rptr_gray[7]_net_1\, rptr_gray(6) => 
        \rptr_gray[6]_net_1\, rptr_gray(5) => 
        \rptr_gray[5]_net_1\, rptr_gray(4) => 
        \rptr_gray[4]_net_1\, rptr_gray(3) => 
        \rptr_gray[3]_net_1\, rptr_gray(2) => 
        \rptr_gray[2]_net_1\, rptr_gray(1) => 
        \rptr_gray[1]_net_1\, rptr_gray(0) => 
        \rptr_gray[0]_net_1\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\, rptr_bin_sync_0 => 
        \rptr_bin_sync[11]\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, itx_fifo_rst_i => 
        itx_fifo_rst_i);
    
    wptr_s_267 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => wptr_s_267_FCO);
    
    \rptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[3]_net_1\, S
         => \rptr_s[4]\, Y => OPEN, FCO => \rptr_cry[4]_net_1\);
    
    wdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[2]_net_1\, B => 
        \rptr_bin_sync2[2]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_1\, S => \wdiff_bus[2]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_2\);
    
    \rptr_gray[2]\ : SLE
      port map(D => \rptr_gray_1[2]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[2]_net_1\);
    
    \wptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[8]_net_1\, S
         => \wptr_s[9]\, Y => OPEN, FCO => \wptr_cry[9]_net_1\);
    
    \wptr_bin_sync2[3]\ : SLE
      port map(D => \wptr_bin_sync[3]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[3]_net_1\);
    
    \wptr[2]\ : SLE
      port map(D => \wptr_s[2]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[2]_net_1\);
    
    \rptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[1]_net_1\, S
         => \rptr_s[2]\, Y => OPEN, FCO => \rptr_cry[2]_net_1\);
    
    rdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[9]_net_1\, B => 
        \rptr[9]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_8\, S => \rdiff_bus[9]\, Y => OPEN, FCO
         => \rdiff_bus_cry_9\);
    
    \memwaddr_r[0]\ : SLE
      port map(D => \memwaddr_r_s[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[0]\);
    
    \wptr_gray[2]\ : SLE
      port map(D => \wptr_gray_1[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[2]_net_1\);
    
    wdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[4]_net_1\, B => 
        \rptr_bin_sync2[4]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_3\, S => \wdiff_bus[4]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_4\);
    
    \memwaddr_r_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[1]_net_1\, S => \memwaddr_r_s[2]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[2]_net_1\);
    
    \wptr_gray[11]\ : SLE
      port map(D => \wptr[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[9]\ : SLE
      port map(D => \wptr_bin_sync[9]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[9]_net_1\);
    
    \rptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[6]_net_1\, B => \rptr[7]_net_1\, Y => 
        \rptr_gray_1[6]_net_1\);
    
    \wptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[11]_net_1\, B => \wptr[10]_net_1\, Y
         => \wptr_gray_1[10]_net_1\);
    
    wdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[6]_net_1\, B => 
        \rptr_bin_sync2[6]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_5\, S => \wdiff_bus[6]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_6\);
    
    memwaddr_r_s_269 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => memwaddr_r_s_269_FCO);
    
    \rptr_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[10]_net_1\, S
         => \rptr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \rptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[2]_net_1\, S
         => \rptr_s[3]\, Y => OPEN, FCO => \rptr_cry[3]_net_1\);
    
    \memraddr_r[4]\ : SLE
      port map(D => \memraddr_r_s[4]\, CLK => BIT_CLK, EN => 
        fifo_MEMRE, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[4]\);
    
    \memraddr_r_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[6]_net_1\, S => \memraddr_r_s[7]\, Y => 
        OPEN, FCO => \memraddr_r_cry[7]_net_1\);
    
    \memraddr_r_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[8]_net_1\, S => \memraddr_r_s[9]\, Y => 
        OPEN, FCO => \memraddr_r_cry[9]_net_1\);
    
    \memraddr_r[5]\ : SLE
      port map(D => \memraddr_r_s[5]\, CLK => BIT_CLK, EN => 
        fifo_MEMRE, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[5]\);
    
    \rptr_gray[6]\ : SLE
      port map(D => \rptr_gray_1[6]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[6]_net_1\);
    
    \memraddr_r[9]\ : SLE
      port map(D => \memraddr_r_s[9]\, CLK => BIT_CLK, EN => 
        fifo_MEMRE, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[9]\);
    
    \rptr[0]\ : SLE
      port map(D => \rptr_s[0]\, CLK => BIT_CLK, EN => fifo_MEMRE, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[0]_net_1\);
    
    \wptr[10]\ : SLE
      port map(D => \wptr_s[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \wptr[10]_net_1\);
    
    \memwaddr_r_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[3]_net_1\, S => \memwaddr_r_s[4]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[4]_net_1\);
    
    \memraddr_r_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[2]_net_1\, S => \memraddr_r_s[3]\, Y => 
        OPEN, FCO => \memraddr_r_cry[3]_net_1\);
    
    wdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[1]_net_1\, B => 
        \rptr_bin_sync2[1]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_0\, S => \wdiff_bus[1]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_1\);
    
    rdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[2]_net_1\, B => 
        \rptr[2]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_1\, S => \rdiff_bus[2]\, Y => OPEN, FCO
         => \rdiff_bus_cry_2\);
    
    \wptr_gray[9]\ : SLE
      port map(D => \wptr_gray_1[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[9]_net_1\);
    
    \rptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[4]_net_1\, B => \rptr[5]_net_1\, Y => 
        \rptr_gray_1[4]_net_1\);
    
    \wptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[8]_net_1\, B => \wptr[9]_net_1\, Y => 
        \wptr_gray_1[8]_net_1\);
    
    Rd_corefifo_grayToBinConv : 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv
      port map(rptr_bin_sync(11) => \rptr_bin_sync[11]\, 
        rptr_bin_sync(10) => \rptr_bin_sync[10]\, 
        rptr_bin_sync(9) => \rptr_bin_sync[9]\, rptr_bin_sync(8)
         => \rptr_bin_sync[8]\, rptr_bin_sync(7) => 
        \rptr_bin_sync[7]\, rptr_bin_sync(6) => 
        \rptr_bin_sync[6]\, rptr_bin_sync(5) => 
        \rptr_bin_sync[5]\, rptr_bin_sync(4) => 
        \rptr_bin_sync[4]\, rptr_bin_sync(3) => 
        \rptr_bin_sync[3]\, rptr_bin_sync(2) => 
        \rptr_bin_sync[2]\, rptr_bin_sync(1) => 
        \rptr_bin_sync[1]\, rptr_bin_sync(0) => 
        \rptr_bin_sync[0]\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\);
    
    \rptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => rptr_s_268_FCO, S => 
        \rptr_s[1]\, Y => OPEN, FCO => \rptr_cry[1]_net_1\);
    
    rdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[3]_net_1\, B => 
        \rptr[3]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_2\, S => \rdiff_bus[3]\, Y => OPEN, FCO
         => \rdiff_bus_cry_3\);
    
    rdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[10]_net_1\, B => 
        \rptr[10]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_9\, S => \rdiff_bus[10]\, Y => OPEN, FCO
         => \rdiff_bus_cry_10\);
    
    \memraddr_r_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[5]_net_1\, S => \memraddr_r_s[6]\, Y => 
        OPEN, FCO => \memraddr_r_cry[6]_net_1\);
    
    \memraddr_r[6]\ : SLE
      port map(D => \memraddr_r_s[6]\, CLK => BIT_CLK, EN => 
        fifo_MEMRE, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[6]\);
    
    \rptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[6]_net_1\, S
         => \rptr_s[7]\, Y => OPEN, FCO => \rptr_cry[7]_net_1\);
    
    rdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => rdiff_bus, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => rdiff_bus_cry_0_Y, FCO => \rdiff_bus_cry_0\);
    
    memraddr_r_s_270 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => memraddr_r_s_270_FCO);
    
    \memraddr_r[2]\ : SLE
      port map(D => \memraddr_r_s[2]\, CLK => BIT_CLK, EN => 
        fifo_MEMRE, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[2]\);
    
    \wptr[8]\ : SLE
      port map(D => \wptr_s[8]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[8]_net_1\);
    
    wdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[3]_net_1\, B => 
        \rptr_bin_sync2[3]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_2\, S => \wdiff_bus[3]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_3\);
    
    \rptr_gray[7]\ : SLE
      port map(D => \rptr_gray_1[7]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[7]_net_1\);
    
    \wptr_gray[0]\ : SLE
      port map(D => \wptr_gray_1[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[0]_net_1\);
    
    \rptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[0]_net_1\, B => \rptr[1]_net_1\, Y => 
        \rptr_gray_1[0]_net_1\);
    
    \rptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[8]_net_1\, B => \rptr[9]_net_1\, Y => 
        \rptr_gray_1[8]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO is

    port( CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          TX_FIFO_UNDERRUN             : out   std_logic;
          TX_FIFO_UNDERRUN_i           : out   std_logic;
          TX_FIFO_OVERFLOW             : out   std_logic;
          TX_FIFO_OVERFLOW_i           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic;
          un2_re_p                     : in    std_logic;
          TX_FIFO_Empty                : out   std_logic;
          TX_FIFO_Full                 : out   std_logic;
          TX_FIFO_wr_en                : in    std_logic;
          N_516                        : out   std_logic;
          N_517                        : out   std_logic;
          N_518                        : out   std_logic;
          N_519                        : out   std_logic;
          N_520                        : out   std_logic;
          N_521                        : out   std_logic;
          N_228                        : out   std_logic;
          N_522                        : out   std_logic;
          TX_FIFO_rd_en                : in    std_logic;
          fifo_MEMRE                   : in    std_logic;
          m34                          : in    std_logic;
          REN_d1                       : out   std_logic;
          m35                          : in    std_logic;
          BIT_CLK                      : in    std_logic;
          itx_fifo_rst_i               : in    std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO;

architecture DEF_ARCH of FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper
    port( RDATA_int                    : out   std_logic_vector(7 downto 0);
          fifo_MEMRADDR                : in    std_logic_vector(10 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          fifo_MEMWADDR                : in    std_logic_vector(10 downto 0) := (others => 'U');
          BIT_CLK                      : in    std_logic := 'U';
          fifo_MEMRE                   : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic := 'U';
          fifo_MEMWE                   : in    std_logic := 'U'
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async
    port( fifo_MEMWADDR             : out   std_logic_vector(10 downto 0);
          fifo_MEMRADDR             : out   std_logic_vector(10 downto 0);
          TX_FIFO_rd_en             : in    std_logic := 'U';
          TX_FIFO_wr_en             : in    std_logic := 'U';
          fifo_MEMWE                : out   std_logic;
          fifo_MEMRE                : in    std_logic := 'U';
          TX_FIFO_Full              : out   std_logic;
          TX_FIFO_Empty             : out   std_logic;
          un2_re_p                  : in    std_logic := 'U';
          BIT_CLK                   : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          itx_fifo_rst_i            : in    std_logic := 'U';
          TX_FIFO_OVERFLOW_i        : out   std_logic;
          TX_FIFO_OVERFLOW          : out   std_logic;
          TX_FIFO_UNDERRUN_i        : out   std_logic;
          TX_FIFO_UNDERRUN          : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \RDATA_r[5]_net_1\, VCC_net_1, \RDATA_int[5]\, 
        GND_net_1, \RDATA_r[6]_net_1\, \RDATA_int[6]\, 
        \RDATA_r[7]_net_1\, \RDATA_int[7]\, \re_set\, 
        REN_d1_net_1, \RDATA_r[0]_net_1\, \RDATA_int[0]\, 
        \RDATA_r[1]_net_1\, \RDATA_int[1]\, \RDATA_r[2]_net_1\, 
        \RDATA_int[2]\, \RDATA_r[3]_net_1\, \RDATA_int[3]\, 
        \RDATA_r[4]_net_1\, \RDATA_int[4]\, \RE_d1\, 
        \re_pulse_d1\, \re_pulse\, \fifo_MEMWADDR[0]\, 
        \fifo_MEMWADDR[1]\, \fifo_MEMWADDR[2]\, 
        \fifo_MEMWADDR[3]\, \fifo_MEMWADDR[4]\, 
        \fifo_MEMWADDR[5]\, \fifo_MEMWADDR[6]\, 
        \fifo_MEMWADDR[7]\, \fifo_MEMWADDR[8]\, 
        \fifo_MEMWADDR[9]\, \fifo_MEMWADDR[10]\, 
        \fifo_MEMRADDR[0]\, \fifo_MEMRADDR[1]\, 
        \fifo_MEMRADDR[2]\, \fifo_MEMRADDR[3]\, 
        \fifo_MEMRADDR[4]\, \fifo_MEMRADDR[5]\, 
        \fifo_MEMRADDR[6]\, \fifo_MEMRADDR[7]\, 
        \fifo_MEMRADDR[8]\, \fifo_MEMRADDR[9]\, 
        \fifo_MEMRADDR[10]\, fifo_MEMWE : std_logic;

    for all : FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper
	Use entity work.FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper(DEF_ARCH);
    for all : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async
	Use entity work.FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async(DEF_ARCH);
begin 

    REN_d1 <= REN_d1_net_1;

    re_pulse : CFG2
      generic map(INIT => x"E")

      port map(A => m35, B => \re_set\, Y => \re_pulse\);
    
    \RDATA_r[3]\ : SLE
      port map(D => \RDATA_int[3]\, CLK => BIT_CLK, EN => m35, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[3]_net_1\);
    
    \Q_i_m2[2]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[2]_net_1\, C => 
        \RDATA_int[2]\, D => \RE_d1\, Y => N_518);
    
    re_pulse_d1 : SLE
      port map(D => \re_pulse\, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \re_pulse_d1\);
    
    \RDATA_r[5]\ : SLE
      port map(D => \RDATA_int[5]\, CLK => BIT_CLK, EN => m35, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[5]_net_1\);
    
    \Q_i_m2[0]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[0]_net_1\, C => 
        \RDATA_int[0]\, D => \RE_d1\, Y => N_516);
    
    \Q_i_m2[3]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[3]_net_1\, C => 
        \RDATA_int[3]\, D => \RE_d1\, Y => N_519);
    
    \Q_i_m2[7]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[7]_net_1\, C => 
        \RDATA_int[7]\, D => \RE_d1\, Y => N_522);
    
    \Q_i_m2[6]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[6]_net_1\, C => 
        \RDATA_int[6]\, D => \RE_d1\, Y => N_228);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \RW1.UI_ram_wrapper_1\ : FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper
      port map(RDATA_int(7) => \RDATA_int[7]\, RDATA_int(6) => 
        \RDATA_int[6]\, RDATA_int(5) => \RDATA_int[5]\, 
        RDATA_int(4) => \RDATA_int[4]\, RDATA_int(3) => 
        \RDATA_int[3]\, RDATA_int(2) => \RDATA_int[2]\, 
        RDATA_int(1) => \RDATA_int[1]\, RDATA_int(0) => 
        \RDATA_int[0]\, fifo_MEMRADDR(10) => \fifo_MEMRADDR[10]\, 
        fifo_MEMRADDR(9) => \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8)
         => \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), fifo_MEMWADDR(10) => 
        \fifo_MEMWADDR[10]\, fifo_MEMWADDR(9) => 
        \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8) => 
        \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, BIT_CLK => BIT_CLK, fifo_MEMRE => 
        fifo_MEMRE, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, fifo_MEMWE => fifo_MEMWE);
    
    \RDATA_r[0]\ : SLE
      port map(D => \RDATA_int[0]\, CLK => BIT_CLK, EN => m35, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[0]_net_1\);
    
    \Q_i_m2[5]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[5]_net_1\, C => 
        \RDATA_int[5]\, D => \RE_d1\, Y => N_521);
    
    \RDATA_r[2]\ : SLE
      port map(D => \RDATA_int[2]\, CLK => BIT_CLK, EN => m35, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[2]_net_1\);
    
    \Q_i_m2[1]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[1]_net_1\, C => 
        \RDATA_int[1]\, D => \RE_d1\, Y => N_517);
    
    \RDATA_r[6]\ : SLE
      port map(D => \RDATA_int[6]\, CLK => BIT_CLK, EN => m35, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[6]_net_1\);
    
    \L31.U_corefifo_async\ : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async
      port map(fifo_MEMWADDR(10) => \fifo_MEMWADDR[10]\, 
        fifo_MEMWADDR(9) => \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8)
         => \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, fifo_MEMRADDR(10) => 
        \fifo_MEMRADDR[10]\, fifo_MEMRADDR(9) => 
        \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8) => 
        \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, TX_FIFO_rd_en => TX_FIFO_rd_en, 
        TX_FIFO_wr_en => TX_FIFO_wr_en, fifo_MEMWE => fifo_MEMWE, 
        fifo_MEMRE => fifo_MEMRE, TX_FIFO_Full => TX_FIFO_Full, 
        TX_FIFO_Empty => TX_FIFO_Empty, un2_re_p => un2_re_p, 
        BIT_CLK => BIT_CLK, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, itx_fifo_rst_i => 
        itx_fifo_rst_i, TX_FIFO_OVERFLOW_i => TX_FIFO_OVERFLOW_i, 
        TX_FIFO_OVERFLOW => TX_FIFO_OVERFLOW, TX_FIFO_UNDERRUN_i
         => TX_FIFO_UNDERRUN_i, TX_FIFO_UNDERRUN => 
        TX_FIFO_UNDERRUN);
    
    re_set : SLE
      port map(D => REN_d1_net_1, CLK => BIT_CLK, EN => m34, ALn
         => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \re_set\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    RE_d1 : SLE
      port map(D => TX_FIFO_rd_en, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RE_d1\);
    
    \RDATA_r[7]\ : SLE
      port map(D => \RDATA_int[7]\, CLK => BIT_CLK, EN => m35, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[7]_net_1\);
    
    \RDATA_r[4]\ : SLE
      port map(D => \RDATA_int[4]\, CLK => BIT_CLK, EN => m35, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[4]_net_1\);
    
    \REN_d1\ : SLE
      port map(D => fifo_MEMRE, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => REN_d1_net_1);
    
    \Q_i_m2[4]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[4]_net_1\, C => 
        \RDATA_int[4]\, D => \RE_d1\, Y => N_520);
    
    \RDATA_r[1]\ : SLE
      port map(D => \RDATA_int[1]\, CLK => BIT_CLK, EN => m35, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[1]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8 is

    port( CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          itx_fifo_rst_i               : in    std_logic;
          BIT_CLK                      : in    std_logic;
          m35                          : in    std_logic;
          REN_d1                       : out   std_logic;
          m34                          : in    std_logic;
          fifo_MEMRE                   : in    std_logic;
          TX_FIFO_rd_en                : in    std_logic;
          N_522                        : out   std_logic;
          N_228                        : out   std_logic;
          N_521                        : out   std_logic;
          N_520                        : out   std_logic;
          N_519                        : out   std_logic;
          N_518                        : out   std_logic;
          N_517                        : out   std_logic;
          N_516                        : out   std_logic;
          TX_FIFO_wr_en                : in    std_logic;
          TX_FIFO_Full                 : out   std_logic;
          TX_FIFO_Empty                : out   std_logic;
          un2_re_p                     : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic;
          TX_FIFO_OVERFLOW_i           : out   std_logic;
          TX_FIFO_OVERFLOW             : out   std_logic;
          TX_FIFO_UNDERRUN_i           : out   std_logic;
          TX_FIFO_UNDERRUN             : out   std_logic
        );

end FIFO_2Kx8;

architecture DEF_ARCH of FIFO_2Kx8 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO
    port( CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          TX_FIFO_UNDERRUN             : out   std_logic;
          TX_FIFO_UNDERRUN_i           : out   std_logic;
          TX_FIFO_OVERFLOW             : out   std_logic;
          TX_FIFO_OVERFLOW_i           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic := 'U';
          un2_re_p                     : in    std_logic := 'U';
          TX_FIFO_Empty                : out   std_logic;
          TX_FIFO_Full                 : out   std_logic;
          TX_FIFO_wr_en                : in    std_logic := 'U';
          N_516                        : out   std_logic;
          N_517                        : out   std_logic;
          N_518                        : out   std_logic;
          N_519                        : out   std_logic;
          N_520                        : out   std_logic;
          N_521                        : out   std_logic;
          N_228                        : out   std_logic;
          N_522                        : out   std_logic;
          TX_FIFO_rd_en                : in    std_logic := 'U';
          fifo_MEMRE                   : in    std_logic := 'U';
          m34                          : in    std_logic := 'U';
          REN_d1                       : out   std_logic;
          m35                          : in    std_logic := 'U';
          BIT_CLK                      : in    std_logic := 'U';
          itx_fifo_rst_i               : in    std_logic := 'U'
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO
	Use entity work.FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    FIFO_2Kx8_0 : FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO
      port map(CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), TX_FIFO_UNDERRUN => 
        TX_FIFO_UNDERRUN, TX_FIFO_UNDERRUN_i => 
        TX_FIFO_UNDERRUN_i, TX_FIFO_OVERFLOW => TX_FIFO_OVERFLOW, 
        TX_FIFO_OVERFLOW_i => TX_FIFO_OVERFLOW_i, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        un2_re_p => un2_re_p, TX_FIFO_Empty => TX_FIFO_Empty, 
        TX_FIFO_Full => TX_FIFO_Full, TX_FIFO_wr_en => 
        TX_FIFO_wr_en, N_516 => N_516, N_517 => N_517, N_518 => 
        N_518, N_519 => N_519, N_520 => N_520, N_521 => N_521, 
        N_228 => N_228, N_522 => N_522, TX_FIFO_rd_en => 
        TX_FIFO_rd_en, fifo_MEMRE => fifo_MEMRE, m34 => m34, 
        REN_d1 => REN_d1, m35 => m35, BIT_CLK => BIT_CLK, 
        itx_fifo_rst_i => itx_fifo_rst_i);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFOs is

    port( RX_FIFO_DIN_pipe             : in    std_logic_vector(8 downto 0);
          rdiff_bus                    : out   std_logic_vector(13 downto 1);
          RDATA_int                    : out   std_logic_vector(7 downto 0);
          RDATA_r                      : out   std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          RX_FIFO_UNDERRUN             : out   std_logic;
          RX_FIFO_UNDERRUN_i           : out   std_logic;
          RX_FIFO_OVERFLOW             : out   std_logic;
          RX_FIFO_OVERFLOW_i           : out   std_logic;
          CommsFPGA_CCC_0_GL0          : in    std_logic;
          RX_FIFO_Empty                : out   std_logic;
          empty_r_3                    : in    std_logic;
          RX_FIFO_Full                 : out   std_logic;
          un2_re_p_0                   : in    std_logic;
          rdiff_bus_cry_0_Y_0          : out   std_logic;
          iRX_FIFO_wr_en               : in    std_logic;
          sampler_clk1x_en             : in    std_logic;
          RX_InProcess_d1              : in    std_logic;
          tx_col_detect_en             : in    std_logic;
          N_357                        : out   std_logic;
          re_pulse_d1                  : out   std_logic;
          RX_FIFO_rd_en                : in    std_logic;
          RE_d1                        : out   std_logic;
          N_283_i                      : in    std_logic;
          N_314_i_i                    : in    std_logic;
          REN_d1_0                     : out   std_logic;
          iRX_FIFO_rd_en_RNIJFNA_0     : in    std_logic;
          TX_FIFO_UNDERRUN             : out   std_logic;
          TX_FIFO_UNDERRUN_i           : out   std_logic;
          TX_FIFO_OVERFLOW             : out   std_logic;
          TX_FIFO_OVERFLOW_i           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic;
          un2_re_p                     : in    std_logic;
          TX_FIFO_Empty                : out   std_logic;
          TX_FIFO_Full                 : out   std_logic;
          TX_FIFO_wr_en                : in    std_logic;
          N_516                        : out   std_logic;
          N_517                        : out   std_logic;
          N_518                        : out   std_logic;
          N_519                        : out   std_logic;
          N_520                        : out   std_logic;
          N_521                        : out   std_logic;
          N_228                        : out   std_logic;
          N_522                        : out   std_logic;
          TX_FIFO_rd_en                : in    std_logic;
          fifo_MEMRE                   : in    std_logic;
          m34                          : in    std_logic;
          REN_d1                       : out   std_logic;
          m35                          : in    std_logic;
          BIT_CLK                      : in    std_logic;
          RX_FIFO_RST                  : in    std_logic;
          TX_FIFO_RST                  : in    std_logic;
          N_480                        : in    std_logic
        );

end FIFOs;

architecture DEF_ARCH of FIFOs is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9
    port( RDATA_r                   : out   std_logic_vector(7 downto 0);
          RDATA_int                 : out   std_logic_vector(7 downto 0);
          rdiff_bus                 : out   std_logic_vector(13 downto 1);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          irx_fifo_rst_i            : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          iRX_FIFO_rd_en_RNIJFNA_0  : in    std_logic := 'U';
          REN_d1                    : out   std_logic;
          N_314_i_i                 : in    std_logic := 'U';
          N_283_i                   : in    std_logic := 'U';
          RE_d1                     : out   std_logic;
          RX_FIFO_rd_en             : in    std_logic := 'U';
          re_pulse_d1               : out   std_logic;
          N_357                     : out   std_logic;
          tx_col_detect_en          : in    std_logic := 'U';
          RX_InProcess_d1           : in    std_logic := 'U';
          sampler_clk1x_en          : in    std_logic := 'U';
          iRX_FIFO_wr_en            : in    std_logic := 'U';
          rdiff_bus_cry_0_Y_0       : out   std_logic;
          un2_re_p                  : in    std_logic := 'U';
          RX_FIFO_Full              : out   std_logic;
          empty_r_3                 : in    std_logic := 'U';
          RX_FIFO_Empty             : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          RX_FIFO_OVERFLOW_i        : out   std_logic;
          RX_FIFO_OVERFLOW          : out   std_logic;
          RX_FIFO_UNDERRUN_i        : out   std_logic;
          RX_FIFO_UNDERRUN          : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8
    port( CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          itx_fifo_rst_i               : in    std_logic := 'U';
          BIT_CLK                      : in    std_logic := 'U';
          m35                          : in    std_logic := 'U';
          REN_d1                       : out   std_logic;
          m34                          : in    std_logic := 'U';
          fifo_MEMRE                   : in    std_logic := 'U';
          TX_FIFO_rd_en                : in    std_logic := 'U';
          N_522                        : out   std_logic;
          N_228                        : out   std_logic;
          N_521                        : out   std_logic;
          N_520                        : out   std_logic;
          N_519                        : out   std_logic;
          N_518                        : out   std_logic;
          N_517                        : out   std_logic;
          N_516                        : out   std_logic;
          TX_FIFO_wr_en                : in    std_logic := 'U';
          TX_FIFO_Full                 : out   std_logic;
          TX_FIFO_Empty                : out   std_logic;
          un2_re_p                     : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic := 'U';
          TX_FIFO_OVERFLOW_i           : out   std_logic;
          TX_FIFO_OVERFLOW             : out   std_logic;
          TX_FIFO_UNDERRUN_i           : out   std_logic;
          TX_FIFO_UNDERRUN             : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal itx_fifo_rst_i, \itx_fifo_rst\, irx_fifo_rst_i, 
        \irx_fifo_rst\, GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9
	Use entity work.FIFO_8Kx9(DEF_ARCH);
    for all : FIFO_2Kx8
	Use entity work.FIFO_2Kx8(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    irx_fifo_rst : CFG2
      generic map(INIT => x"1")

      port map(A => N_480, B => RX_FIFO_RST, Y => \irx_fifo_rst\);
    
    RECEIVE_FIFO : FIFO_8Kx9
      port map(RDATA_r(7) => RDATA_r(7), RDATA_r(6) => RDATA_r(6), 
        RDATA_r(5) => RDATA_r(5), RDATA_r(4) => RDATA_r(4), 
        RDATA_r(3) => RDATA_r(3), RDATA_r(2) => RDATA_r(2), 
        RDATA_r(1) => RDATA_r(1), RDATA_r(0) => RDATA_r(0), 
        RDATA_int(7) => RDATA_int(7), RDATA_int(6) => 
        RDATA_int(6), RDATA_int(5) => RDATA_int(5), RDATA_int(4)
         => RDATA_int(4), RDATA_int(3) => RDATA_int(3), 
        RDATA_int(2) => RDATA_int(2), RDATA_int(1) => 
        RDATA_int(1), RDATA_int(0) => RDATA_int(0), rdiff_bus(13)
         => rdiff_bus(13), rdiff_bus(12) => rdiff_bus(12), 
        rdiff_bus(11) => rdiff_bus(11), rdiff_bus(10) => 
        rdiff_bus(10), rdiff_bus(9) => rdiff_bus(9), rdiff_bus(8)
         => rdiff_bus(8), rdiff_bus(7) => rdiff_bus(7), 
        rdiff_bus(6) => rdiff_bus(6), rdiff_bus(5) => 
        rdiff_bus(5), rdiff_bus(4) => rdiff_bus(4), rdiff_bus(3)
         => rdiff_bus(3), rdiff_bus(2) => rdiff_bus(2), 
        rdiff_bus(1) => rdiff_bus(1), RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), irx_fifo_rst_i => irx_fifo_rst_i, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        iRX_FIFO_rd_en_RNIJFNA_0 => iRX_FIFO_rd_en_RNIJFNA_0, 
        REN_d1 => REN_d1_0, N_314_i_i => N_314_i_i, N_283_i => 
        N_283_i, RE_d1 => RE_d1, RX_FIFO_rd_en => RX_FIFO_rd_en, 
        re_pulse_d1 => re_pulse_d1, N_357 => N_357, 
        tx_col_detect_en => tx_col_detect_en, RX_InProcess_d1 => 
        RX_InProcess_d1, sampler_clk1x_en => sampler_clk1x_en, 
        iRX_FIFO_wr_en => iRX_FIFO_wr_en, rdiff_bus_cry_0_Y_0 => 
        rdiff_bus_cry_0_Y_0, un2_re_p => un2_re_p_0, RX_FIFO_Full
         => RX_FIFO_Full, empty_r_3 => empty_r_3, RX_FIFO_Empty
         => RX_FIFO_Empty, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, RX_FIFO_OVERFLOW_i => 
        RX_FIFO_OVERFLOW_i, RX_FIFO_OVERFLOW => RX_FIFO_OVERFLOW, 
        RX_FIFO_UNDERRUN_i => RX_FIFO_UNDERRUN_i, 
        RX_FIFO_UNDERRUN => RX_FIFO_UNDERRUN);
    
    itx_fifo_rst : CFG2
      generic map(INIT => x"1")

      port map(A => N_480, B => TX_FIFO_RST, Y => \itx_fifo_rst\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    TRANSMIT_FIFO : FIFO_2Kx8
      port map(CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), itx_fifo_rst_i => 
        itx_fifo_rst_i, BIT_CLK => BIT_CLK, m35 => m35, REN_d1
         => REN_d1, m34 => m34, fifo_MEMRE => fifo_MEMRE, 
        TX_FIFO_rd_en => TX_FIFO_rd_en, N_522 => N_522, N_228 => 
        N_228, N_521 => N_521, N_520 => N_520, N_519 => N_519, 
        N_518 => N_518, N_517 => N_517, N_516 => N_516, 
        TX_FIFO_wr_en => TX_FIFO_wr_en, TX_FIFO_Full => 
        TX_FIFO_Full, TX_FIFO_Empty => TX_FIFO_Empty, un2_re_p
         => un2_re_p, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, TX_FIFO_OVERFLOW_i => 
        TX_FIFO_OVERFLOW_i, TX_FIFO_OVERFLOW => TX_FIFO_OVERFLOW, 
        TX_FIFO_UNDERRUN_i => TX_FIFO_UNDERRUN_i, 
        TX_FIFO_UNDERRUN => TX_FIFO_UNDERRUN);
    
    itx_fifo_rst_RNIUMSA : CLKINT
      port map(A => \itx_fifo_rst\, Y => itx_fifo_rst_i);
    
    irx_fifo_rst_RNIS228 : CLKINT
      port map(A => \irx_fifo_rst\, Y => irx_fifo_rst_i);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Interrupts is

    port( CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PADDR  : in    std_logic_vector(5 downto 2);
          i_int_mask_reg               : in    std_logic_vector(7 downto 0);
          int_reg_6                    : out   std_logic;
          int_reg_3                    : out   std_logic;
          int_reg_0                    : out   std_logic;
          int_reg_4                    : out   std_logic;
          N_26                         : in    std_logic;
          CommsFPGA_top_0_INT          : out   std_logic;
          N_238                        : out   std_logic;
          long_reset                   : in    std_logic;
          CommsFPGA_CCC_0_LOCK         : in    std_logic;
          write_reg_en                 : in    std_logic;
          un29_int_reg_clr             : out   std_logic;
          N_480_rs                     : in    std_logic;
          rx_CRC_error_set             : in    std_logic;
          un33_int_reg_clr             : out   std_logic;
          col_detect_int               : out   std_logic;
          N_480_rs_0                   : in    std_logic;
          TX_collision_detect_set      : in    std_logic;
          rx_packet_complt             : in    std_logic;
          un9_int_reg_clr              : out   std_logic;
          rx_packet_avail_int          : out   std_logic;
          rx_packet_complt_set         : in    std_logic;
          un13_int_reg_clr             : out   std_logic;
          N_480_rs_1                   : in    std_logic;
          TX_FIFO_UNDERRUN_set         : in    std_logic;
          un17_int_reg_clr             : out   std_logic;
          N_480_rs_2                   : in    std_logic;
          TX_FIFO_OVERFLOW_set         : in    std_logic;
          un21_int_reg_clr             : out   std_logic;
          rx_FIFO_UNDERRUN_int         : out   std_logic;
          N_480_rs_3                   : in    std_logic;
          RX_FIFO_UNDERRUN_set         : in    std_logic;
          un25_int_reg_clr             : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic;
          rx_FIFO_OVERFLOW_int         : out   std_logic;
          N_480_rs_4                   : in    std_logic;
          RX_FIFO_OVERFLOW_set         : in    std_logic;
          tx_packet_complt             : in    std_logic;
          CommsFPGA_CCC_0_GL0          : in    std_logic;
          N_480_i                      : out   std_logic;
          N_480                        : out   std_logic;
          N_9_0_i_i                    : out   std_logic
        );

end Interrupts;

architecture DEF_ARCH of Interrupts is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \RESET_i_a2_RNIC0QJ\, \N_480\, \RESET_i_a2\, 
        \N_480_i\, \tx_packet_complt_toClk16x\, 
        tx_packet_complt_toClk16x_i, 
        \tx_packet_complt_d[0]_net_1\, VCC_net_1, GND_net_1, 
        \tx_packet_complt_d[1]_net_1\, 
        \tx_packet_complt_d[2]_net_1\, 
        \tx_packet_complt_d[3]_net_1\, 
        \tx_packet_complt_d[4]_net_1\, 
        \tx_packet_complt_d[5]_net_1\, 
        \tx_packet_complt_d[6]_net_1\, 
        \tx_packet_complt_d[7]_net_1\, rx_FIFO_OVERFLOW_intrs, 
        rx_FIFO_OVERFLOW_int_net_1, \un25_int_reg_clr\, 
        rx_FIFO_UNDERRUN_intrs, rx_FIFO_UNDERRUN_int_net_1, 
        \un21_int_reg_clr\, tx_FIFO_OVERFLOW_intrs, 
        \tx_FIFO_OVERFLOW_int\, \un17_int_reg_clr\, 
        tx_FIFO_UNDERRUN_intrs, \tx_FIFO_UNDERRUN_int\, 
        \un13_int_reg_clr\, rx_packet_avail_intrs, 
        un15_apb3_reset_rs, rx_packet_avail_int_net_1, 
        un15_apb3_reset_i, \un9_int_reg_clr\, 
        \tx_packet_complt_toClk16x_set\, tx_packet_complt_intrs, 
        un6_apb3_reset_rs, \tx_packet_complt_int\, 
        un6_apb3_reset_i, un5_int_reg_clr, col_detect_intrs, 
        col_detect_int_net_1, \un33_int_reg_clr\, 
        rx_CRC_error_intrs, \rx_CRC_error_int\, 
        \un29_int_reg_clr\, un13_int_reg_clr_0_a2_0, 
        un33_int_reg_clr_0, \int_reg_6\, \int_reg_3\, \int_reg_0\, 
        \int_reg_4\, \INT_3\, \INT_0\, \N_238\, 
        un1_write_reg_en_0_a2_0, \INT_5\ : std_logic;

begin 

    int_reg_6 <= \int_reg_6\;
    int_reg_3 <= \int_reg_3\;
    int_reg_0 <= \int_reg_0\;
    int_reg_4 <= \int_reg_4\;
    N_238 <= \N_238\;
    un29_int_reg_clr <= \un29_int_reg_clr\;
    un33_int_reg_clr <= \un33_int_reg_clr\;
    col_detect_int <= col_detect_int_net_1;
    un9_int_reg_clr <= \un9_int_reg_clr\;
    rx_packet_avail_int <= rx_packet_avail_int_net_1;
    un13_int_reg_clr <= \un13_int_reg_clr\;
    un17_int_reg_clr <= \un17_int_reg_clr\;
    un21_int_reg_clr <= \un21_int_reg_clr\;
    rx_FIFO_UNDERRUN_int <= rx_FIFO_UNDERRUN_int_net_1;
    un25_int_reg_clr <= \un25_int_reg_clr\;
    rx_FIFO_OVERFLOW_int <= rx_FIFO_OVERFLOW_int_net_1;
    N_480_i <= \N_480_i\;
    N_480 <= \N_480\;

    col_detect_int_RNID9FJ : CFG3
      generic map(INIT => x"EC")

      port map(A => TX_collision_detect_set, B => 
        col_detect_intrs, C => N_480_rs_0, Y => 
        col_detect_int_net_1);
    
    \COLLISION_DETECTION_INTR.un33_int_reg_clr_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(0), B => 
        write_reg_en, Y => un33_int_reg_clr_0);
    
    tx_packet_complt_toClk16x_set_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \tx_packet_complt_toClk16x\, Y => 
        tx_packet_complt_toClk16x_i);
    
    \RX_FIFO_UNDERRUN_INTR.un21_int_reg_clr\ : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PWDATA(3), C => 
        un1_write_reg_en_0_a2_0, D => N_26, Y => 
        \un21_int_reg_clr\);
    
    INT_5 : CFG4
      generic map(INIT => x"FFBA")

      port map(A => \int_reg_0\, B => i_int_mask_reg(0), C => 
        col_detect_int_net_1, D => \INT_3\, Y => \INT_5\);
    
    \RX_PACKET_AVAILABLE_INTR.un15_apb3_reset\ : CFG4
      generic map(INIT => x"0001")

      port map(A => rx_FIFO_UNDERRUN_int_net_1, B => 
        rx_FIFO_OVERFLOW_int_net_1, C => \rx_CRC_error_int\, D
         => \N_480\, Y => un15_apb3_reset_i);
    
    \TX_FIFO_UNDERRUN_INTR.un13_int_reg_clr_0_a2_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(5), B => 
        write_reg_en, Y => un13_int_reg_clr_0_a2_0);
    
    \TX_FIFO_OVERFLOW_INTR.un17_int_reg_clr\ : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PWDATA(4), C => 
        un1_write_reg_en_0_a2_0, D => N_26, Y => 
        \un17_int_reg_clr\);
    
    \RX_CRC_ERROR_INTR.un29_int_reg_clr\ : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PWDATA(1), C => 
        un1_write_reg_en_0_a2_0, D => N_26, Y => 
        \un29_int_reg_clr\);
    
    \int_reg_1_RNO[4]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => TX_FIFO_OVERFLOW_set, B => 
        tx_FIFO_OVERFLOW_intrs, C => N_480_rs_2, Y => 
        \tx_FIFO_OVERFLOW_int\);
    
    rx_FIFO_UNDERRUN_int_RNI9TLR : CFG3
      generic map(INIT => x"EC")

      port map(A => RX_FIFO_UNDERRUN_set, B => 
        rx_FIFO_UNDERRUN_intrs, C => N_480_rs_3, Y => 
        rx_FIFO_UNDERRUN_int_net_1);
    
    rx_CRC_error_int_RNIDSP31 : CFG3
      generic map(INIT => x"EC")

      port map(A => rx_CRC_error_set, B => rx_CRC_error_intrs, C
         => N_480_rs, Y => \rx_CRC_error_int\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \rx_packet_avail_int\ : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un9_int_reg_clr\, ALn => un15_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rx_packet_avail_intrs);
    
    \int_reg_1_0_a2_RNO[7]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \tx_packet_complt_toClk16x_set\, B => 
        tx_packet_complt_intrs, C => un6_apb3_reset_rs, Y => 
        \tx_packet_complt_int\);
    
    \tx_packet_complt_d[0]\ : SLE
      port map(D => tx_packet_complt, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => \N_480_i\, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_packet_complt_d[0]_net_1\);
    
    \TX_PACKET_COMPLETE_INTR.un5_int_reg_clr\ : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PWDATA(7), C => 
        un1_write_reg_en_0_a2_0, D => N_26, Y => un5_int_reg_clr);
    
    \tx_packet_complt_d[7]\ : SLE
      port map(D => \tx_packet_complt_d[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => \N_480_i\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_complt_d[7]_net_1\);
    
    tx_FIFO_OVERFLOW_int : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un17_int_reg_clr\, ALn => \N_480_i\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => tx_FIFO_OVERFLOW_intrs);
    
    rx_CRC_error_int : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un29_int_reg_clr\, ALn => \N_480_i\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rx_CRC_error_intrs);
    
    RESET_i_a2_RNIC0QJ : CFG2
      generic map(INIT => x"1")

      port map(A => \N_480\, B => tx_packet_complt, Y => 
        \RESET_i_a2_RNIC0QJ\);
    
    tx_FIFO_UNDERRUN_int : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un13_int_reg_clr\, ALn => \N_480_i\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => tx_FIFO_UNDERRUN_intrs);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \tx_packet_complt_d[5]\ : SLE
      port map(D => \tx_packet_complt_d[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => \N_480_i\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_complt_d[5]_net_1\);
    
    \int_reg_1_0_a2[5]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \tx_FIFO_UNDERRUN_int\, B => 
        i_int_mask_reg(5), Y => \int_reg_4\);
    
    \tx_packet_complt_d[4]\ : SLE
      port map(D => \tx_packet_complt_d[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => \N_480_i\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_complt_d[4]_net_1\);
    
    \REGISTER_CLEAR_INST.un1_write_reg_en_0_a2_0\ : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => \N_238\);
    
    \TX_FIFO_UNDERRUN_INTR.un13_int_reg_clr_0_a2\ : CFG4
      generic map(INIT => x"0800")

      port map(A => \N_238\, B => N_26, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        un13_int_reg_clr_0_a2_0, Y => \un13_int_reg_clr\);
    
    RESET_i_a2_RNIC0QJ_0 : CLKINT
      port map(A => \RESET_i_a2_RNIC0QJ\, Y => N_9_0_i_i);
    
    \REGISTER_CLEAR_INST.un1_write_reg_en_0_a2_0_0\ : CFG4
      generic map(INIT => x"0800")

      port map(A => write_reg_en, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => 
        CoreAPB3_0_APBmslave0_PADDR(5), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => 
        un1_write_reg_en_0_a2_0);
    
    \RX_PACKET_AVAILABLE_INTR.un9_int_reg_clr\ : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PWDATA(6), C => 
        un1_write_reg_en_0_a2_0, D => N_26, Y => 
        \un9_int_reg_clr\);
    
    \RX_PACKET_AVAILABLE_INTR.un15_apb3_reset_rs\ : SLE
      port map(D => VCC_net_1, CLK => rx_packet_complt, EN => 
        VCC_net_1, ALn => un15_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q
         => un15_apb3_reset_rs);
    
    INT_0 : CFG3
      generic map(INIT => x"BA")

      port map(A => \int_reg_6\, B => i_int_mask_reg(6), C => 
        rx_packet_avail_int_net_1, Y => \INT_0\);
    
    \tx_packet_complt_d[3]\ : SLE
      port map(D => \tx_packet_complt_d[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => \N_480_i\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_complt_d[3]_net_1\);
    
    RESET_i_a2_RNISH6E_0 : CFG1
      generic map(INIT => "01")

      port map(A => \N_480\, Y => \N_480_i\);
    
    INT_3 : CFG4
      generic map(INIT => x"7350")

      port map(A => i_int_mask_reg(3), B => i_int_mask_reg(2), C
         => rx_FIFO_UNDERRUN_int_net_1, D => 
        rx_FIFO_OVERFLOW_int_net_1, Y => \INT_3\);
    
    tx_FIFO_UNDERRUN_int_RNIB94L : CFG3
      generic map(INIT => x"EC")

      port map(A => TX_FIFO_UNDERRUN_set, B => 
        tx_FIFO_UNDERRUN_intrs, C => N_480_rs_1, Y => 
        \tx_FIFO_UNDERRUN_int\);
    
    tx_packet_complt_int : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un5_int_reg_clr, ALn => un6_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => tx_packet_complt_intrs);
    
    \int_reg_1_0_a2[7]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \tx_packet_complt_int\, B => 
        i_int_mask_reg(7), Y => \int_reg_6\);
    
    \tx_packet_complt_d[6]\ : SLE
      port map(D => \tx_packet_complt_d[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => \N_480_i\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_complt_d[6]_net_1\);
    
    \int_reg_1[1]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \rx_CRC_error_int\, B => i_int_mask_reg(1), Y
         => \int_reg_0\);
    
    tx_packet_complt_toClk16x : CFG2
      generic map(INIT => x"2")

      port map(A => \tx_packet_complt_d[6]_net_1\, B => 
        \tx_packet_complt_d[7]_net_1\, Y => 
        \tx_packet_complt_toClk16x\);
    
    \rx_FIFO_OVERFLOW_int\ : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un25_int_reg_clr\, ALn => \N_480_i\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rx_FIFO_OVERFLOW_intrs);
    
    RESET_i_a2 : CFG2
      generic map(INIT => x"D")

      port map(A => CommsFPGA_CCC_0_LOCK, B => long_reset, Y => 
        \RESET_i_a2\);
    
    RESET_i_a2_RNISH6E : CLKINT
      port map(A => \RESET_i_a2\, Y => \N_480\);
    
    \tx_packet_complt_d[1]\ : SLE
      port map(D => \tx_packet_complt_d[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => \N_480_i\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_complt_d[1]_net_1\);
    
    rx_FIFO_OVERFLOW_int_RNICNQK : CFG3
      generic map(INIT => x"EC")

      port map(A => RX_FIFO_OVERFLOW_set, B => 
        rx_FIFO_OVERFLOW_intrs, C => N_480_rs_4, Y => 
        rx_FIFO_OVERFLOW_int_net_1);
    
    \tx_packet_complt_d[2]\ : SLE
      port map(D => \tx_packet_complt_d[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => \N_480_i\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_complt_d[2]_net_1\);
    
    \TX_PACKET_COMPLETE_INTR.un6_apb3_reset\ : CFG3
      generic map(INIT => x"01")

      port map(A => \tx_FIFO_UNDERRUN_int\, B => 
        col_detect_int_net_1, C => \N_480\, Y => un6_apb3_reset_i);
    
    \COLLISION_DETECTION_INTR.un33_int_reg_clr\ : CFG4
      generic map(INIT => x"0800")

      port map(A => \N_238\, B => N_26, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => un33_int_reg_clr_0, 
        Y => \un33_int_reg_clr\);
    
    \TX_PACKET_COMPLETE_INTR.un6_apb3_reset_rs\ : SLE
      port map(D => VCC_net_1, CLK => \tx_packet_complt_toClk16x\, 
        EN => VCC_net_1, ALn => un6_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        VCC_net_1, Q => un6_apb3_reset_rs);
    
    INT : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \int_reg_4\, B => \int_reg_3\, C => \INT_5\, 
        D => \INT_0\, Y => CommsFPGA_top_0_INT);
    
    \RX_PACKET_AVAILABLE_INTR.un15_apb3_reset_rs_RNIQI861\ : CFG3
      generic map(INIT => x"EC")

      port map(A => rx_packet_complt_set, B => 
        rx_packet_avail_intrs, C => un15_apb3_reset_rs, Y => 
        rx_packet_avail_int_net_1);
    
    tx_packet_complt_toClk16x_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un5_int_reg_clr, ALn => tx_packet_complt_toClk16x_i, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_complt_toClk16x_set\);
    
    \RX_FIFO_OVERFLOW_INTR.un25_int_reg_clr\ : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PWDATA(2), C => 
        un1_write_reg_en_0_a2_0, D => N_26, Y => 
        \un25_int_reg_clr\);
    
    \int_reg_1[4]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \tx_FIFO_OVERFLOW_int\, B => 
        i_int_mask_reg(4), Y => \int_reg_3\);
    
    \rx_FIFO_UNDERRUN_int\ : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un21_int_reg_clr\, ALn => \N_480_i\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rx_FIFO_UNDERRUN_intrs);
    
    \col_detect_int\ : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un33_int_reg_clr\, ALn => \N_480_i\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => col_detect_intrs);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity uP_if is

    port( rdiff_bus                      : in    std_logic_vector(13 downto 1);
          CoreAPB3_0_APBmslave0_PADDR    : in    std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA_m : out   std_logic_vector(7 downto 0);
          RDATA_int                      : in    std_logic_vector(7 downto 0);
          RDATA_r                        : in    std_logic_vector(7 downto 0);
          consumer_type2_reg             : out   std_logic_vector(9 downto 0);
          consumer_type3_reg             : out   std_logic_vector(9 downto 0);
          consumer_type1_reg             : out   std_logic_vector(9 downto 0);
          consumer_type4_reg             : out   std_logic_vector(9 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA   : in    std_logic_vector(7 downto 0);
          p2s_data_0                     : in    std_logic;
          N_9_0_i_i                      : out   std_logic;
          N_480_i                        : out   std_logic;
          RX_FIFO_OVERFLOW_set           : in    std_logic;
          N_480_rs_4                     : in    std_logic;
          un25_int_reg_clr               : out   std_logic;
          RX_FIFO_UNDERRUN_set           : in    std_logic;
          N_480_rs_3                     : in    std_logic;
          un21_int_reg_clr               : out   std_logic;
          TX_FIFO_OVERFLOW_set           : in    std_logic;
          N_480_rs_2                     : in    std_logic;
          un17_int_reg_clr               : out   std_logic;
          TX_FIFO_UNDERRUN_set           : in    std_logic;
          N_480_rs_1                     : in    std_logic;
          un13_int_reg_clr               : out   std_logic;
          rx_packet_complt_set           : in    std_logic;
          un9_int_reg_clr                : out   std_logic;
          TX_collision_detect_set        : in    std_logic;
          N_480_rs_0                     : in    std_logic;
          un33_int_reg_clr               : out   std_logic;
          rx_CRC_error_set               : in    std_logic;
          N_480_rs                       : in    std_logic;
          un29_int_reg_clr               : out   std_logic;
          CommsFPGA_CCC_0_LOCK           : in    std_logic;
          CommsFPGA_top_0_INT            : out   std_logic;
          empty_r_3                      : out   std_logic;
          N_357                          : in    std_logic;
          tx_packet_complt               : in    std_logic;
          DRVR_EN_c                      : in    std_logic;
          N_209_i                        : out   std_logic;
          rdiff_bus_cry_0_Y_0            : in    std_logic;
          N_314_i_i                      : out   std_logic;
          m34                            : out   std_logic;
          un2_re_p_0                     : out   std_logic;
          TX_FIFO_rd_en                  : in    std_logic;
          CoreAPB3_0_APBmslave0_PENABLE  : in    std_logic;
          CoreAPB3_0_APBmslave0_PWRITE   : in    std_logic;
          iRX_FIFO_rd_en_RNIJFNA_0       : out   std_logic;
          REN_d1_0                       : in    std_logic;
          N_283_i                        : out   std_logic;
          N_6_0                          : out   std_logic;
          N_480                          : out   std_logic;
          TX_PostAmble_d1                : in    std_logic;
          RX_FIFO_RST_1                  : out   std_logic;
          RX_EarlyTerm                   : in    std_logic;
          CoreAPB3_0_APBmslave0_PSELx    : in    std_logic;
          un2_re_p                       : out   std_logic;
          RX_FIFO_Empty                  : in    std_logic;
          TX_FIFO_Full                   : in    std_logic;
          RE_d1                          : in    std_logic;
          re_pulse_d1                    : in    std_logic;
          un19_tx_dataen                 : in    std_logic;
          tx_preamble_pat_en             : in    std_logic;
          TX_PreAmble                    : in    std_logic;
          MANCHESTER_OUT_5               : out   std_logic;
          BIT_CLK                        : in    std_logic;
          fifo_MEMRE                     : out   std_logic;
          m35                            : out   std_logic;
          byte_clk_en                    : in    std_logic;
          REN_d1                         : in    std_logic;
          TX_FIFO_Empty                  : in    std_logic;
          iTX_FIFO_rd_en                 : in    std_logic;
          RX_FIFO_Full                   : in    std_logic;
          rx_packet_complt               : in    std_logic;
          N_386_i_set                    : in    std_logic;
          un25_read_reg_en               : out   std_logic;
          N_386_i_rs                     : in    std_logic;
          TX_FIFO_wr_en                  : out   std_logic;
          N_209_i_i                      : in    std_logic;
          RX_FIFO_rd_en                  : out   std_logic;
          TX_FIFO_RST                    : out   std_logic;
          start_tx_FIFO                  : out   std_logic;
          internal_loopback              : out   std_logic;
          long_reset                     : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY   : out   std_logic;
          long_reset_set                 : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz      : in    std_logic;
          CommsFPGA_CCC_0_GL0            : in    std_logic;
          long_reset_i                   : in    std_logic;
          un2_apb3_addr_13               : out   std_logic;
          N_386_i_i                      : out   std_logic;
          N_106_mux_i_i                  : out   std_logic
        );

end uP_if;

architecture DEF_ARCH of uP_if is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component Interrupts
    port( CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PADDR  : in    std_logic_vector(5 downto 2) := (others => 'U');
          i_int_mask_reg               : in    std_logic_vector(7 downto 0) := (others => 'U');
          int_reg_6                    : out   std_logic;
          int_reg_3                    : out   std_logic;
          int_reg_0                    : out   std_logic;
          int_reg_4                    : out   std_logic;
          N_26                         : in    std_logic := 'U';
          CommsFPGA_top_0_INT          : out   std_logic;
          N_238                        : out   std_logic;
          long_reset                   : in    std_logic := 'U';
          CommsFPGA_CCC_0_LOCK         : in    std_logic := 'U';
          write_reg_en                 : in    std_logic := 'U';
          un29_int_reg_clr             : out   std_logic;
          N_480_rs                     : in    std_logic := 'U';
          rx_CRC_error_set             : in    std_logic := 'U';
          un33_int_reg_clr             : out   std_logic;
          col_detect_int               : out   std_logic;
          N_480_rs_0                   : in    std_logic := 'U';
          TX_collision_detect_set      : in    std_logic := 'U';
          rx_packet_complt             : in    std_logic := 'U';
          un9_int_reg_clr              : out   std_logic;
          rx_packet_avail_int          : out   std_logic;
          rx_packet_complt_set         : in    std_logic := 'U';
          un13_int_reg_clr             : out   std_logic;
          N_480_rs_1                   : in    std_logic := 'U';
          TX_FIFO_UNDERRUN_set         : in    std_logic := 'U';
          un17_int_reg_clr             : out   std_logic;
          N_480_rs_2                   : in    std_logic := 'U';
          TX_FIFO_OVERFLOW_set         : in    std_logic := 'U';
          un21_int_reg_clr             : out   std_logic;
          rx_FIFO_UNDERRUN_int         : out   std_logic;
          N_480_rs_3                   : in    std_logic := 'U';
          RX_FIFO_UNDERRUN_set         : in    std_logic := 'U';
          un25_int_reg_clr             : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic := 'U';
          rx_FIFO_OVERFLOW_int         : out   std_logic;
          N_480_rs_4                   : in    std_logic := 'U';
          RX_FIFO_OVERFLOW_set         : in    std_logic := 'U';
          tx_packet_complt             : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0          : in    std_logic := 'U';
          N_480_i                      : out   std_logic;
          N_480                        : out   std_logic;
          N_9_0_i_i                    : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \control_reg_RNIS9SH1[1]_net_1\, 
        \iAPB3_READY[0]_net_1\, \iAPB3_READY_i[0]\, N_386_i, 
        \N_386_i_i\, un2_apb3_addr_13_net_1, un2_apb3_addr_13_i, 
        \up_EOP_sync[2]_net_1\, VCC_net_1, \up_EOP_sync[1]_net_1\, 
        GND_net_1, \consumer_type3_reg[0]\, 
        un13_address_low3_reg_en, \consumer_type3_reg[1]\, 
        \consumer_type3_reg[2]\, \consumer_type3_reg[3]\, 
        \consumer_type3_reg[4]\, \consumer_type3_reg[5]\, 
        \consumer_type3_reg[6]\, \consumer_type3_reg[7]\, 
        \iAPB3_READYrs[0]\, un5_apb3_rst_rs, un5_apb3_rst_i, 
        CoreAPB3_0_APBmslave0_PREADYrs, 
        \CoreAPB3_0_APBmslave0_PREADY\, \up_EOP_sync[0]_net_1\, 
        \up_EOP\, \consumer_type4_reg[1]\, 
        un13_address_low4_reg_en, \consumer_type4_reg[2]\, 
        \consumer_type4_reg[3]\, \consumer_type4_reg[4]\, 
        \consumer_type4_reg[5]\, \consumer_type4_reg[6]\, 
        \consumer_type4_reg[7]\, \consumer_type4_reg[8]\, 
        un13_address_high4_reg_en, \consumer_type4_reg[9]\, 
        \address_high4_reg[2]_net_1\, 
        \address_high4_reg[3]_net_1\, 
        \address_high4_reg[4]_net_1\, 
        \address_high4_reg[5]_net_1\, 
        \address_high4_reg[6]_net_1\, 
        \address_high4_reg[7]_net_1\, 
        \address_high1_reg[2]_net_1\, un13_address_high1_reg_en, 
        \address_high1_reg[3]_net_1\, 
        \address_high1_reg[4]_net_1\, 
        \address_high1_reg[5]_net_1\, 
        \address_high1_reg[6]_net_1\, 
        \address_high1_reg[7]_net_1\, \control_reg[0]_net_1\, 
        control_reg_105, external_loopback, 
        \control_reg[2]_net_1\, \control_reg[3]_net_1\, 
        \internal_loopback\, \start_tx_FIFO\, N_82_i, 
        un1_control_reg_en_2_i_0, rx_FIFO_rst_reg, \TX_FIFO_RST\, 
        \consumer_type4_reg[0]\, \consumer_type1_reg[3]\, 
        un13_address_low1_reg_en, \consumer_type1_reg[4]\, 
        \consumer_type1_reg[5]\, \consumer_type1_reg[6]\, 
        \consumer_type1_reg[7]\, \scratch_pad_reg[0]_net_1\, 
        \write_scratch_reg_en\, \scratch_pad_reg[1]_net_1\, 
        \scratch_pad_reg[2]_net_1\, \scratch_pad_reg[3]_net_1\, 
        \scratch_pad_reg[4]_net_1\, \scratch_pad_reg[5]_net_1\, 
        \scratch_pad_reg[6]_net_1\, \scratch_pad_reg[7]_net_1\, 
        \consumer_type1_reg[8]\, \consumer_type1_reg[9]\, 
        \consumer_type2_reg[4]\, un13_address_low2_reg_en, 
        \consumer_type2_reg[5]\, \consumer_type2_reg[6]\, 
        \consumer_type2_reg[7]\, \consumer_type2_reg[8]\, 
        un13_address_high2_reg_en, \consumer_type2_reg[9]\, 
        \address_high2_reg[2]_net_1\, 
        \address_high2_reg[3]_net_1\, 
        \address_high2_reg[4]_net_1\, 
        \address_high2_reg[5]_net_1\, 
        \address_high2_reg[6]_net_1\, 
        \address_high2_reg[7]_net_1\, \consumer_type1_reg[0]\, 
        \consumer_type1_reg[1]\, \consumer_type1_reg[2]\, 
        \i_int_mask_reg[5]_net_1\, un13_int_mask_reg_en, 
        \i_int_mask_reg[6]_net_1\, \i_int_mask_reg[7]_net_1\, 
        \consumer_type3_reg[8]\, un13_address_high3_reg_en, 
        \consumer_type3_reg[9]\, \address_high3_reg[2]_net_1\, 
        \address_high3_reg[3]_net_1\, 
        \address_high3_reg[4]_net_1\, 
        \address_high3_reg[5]_net_1\, 
        \address_high3_reg[6]_net_1\, 
        \address_high3_reg[7]_net_1\, \consumer_type2_reg[0]\, 
        \consumer_type2_reg[1]\, \consumer_type2_reg[2]\, 
        \consumer_type2_reg[3]\, \i_int_mask_reg[0]_net_1\, 
        \i_int_mask_reg[1]_net_1\, \i_int_mask_reg[2]_net_1\, 
        \i_int_mask_reg[3]_net_1\, \i_int_mask_reg[4]_net_1\, 
        \RX_FIFO_rd_en\, N_384_i_i, un45_apb3_addr, 
        address_low4_reg_en_1, apb3_addr, \int_mask_reg_en\, 
        un9_apb3_addr, un1_apb3_addr, \control_reg_en\, 
        un5_apb3_addr, \address_low4_reg_en\, un41_apb3_addr, 
        \address_low3_reg_en\, un33_apb3_addr, 
        \address_low2_reg_en\, un25_apb3_addr, 
        \address_low1_reg_en\, un17_apb3_addr, 
        \address_high4_reg_en\, un37_apb3_addr, 
        \address_high3_reg_en\, un29_apb3_addr, 
        \address_high2_reg_en\, un21_apb3_addr, 
        \address_high1_reg_en\, un13_apb3_addr, \write_reg_en\, 
        \read_reg_en\, un53_apb3_addr, \RX_packet_depth_status\, 
        un1_RX_packet_depth_i, \APB3_RDATA_1rs[5]\, 
        \un2_apb3_addr_13_set\, \APB3_RDATA_1[5]_net_1\, 
        \un25_read_reg_en\, \APB3_RDATA_2_i[5]_net_1\, 
        \APB3_RDATA_1rs[6]\, \APB3_RDATA_1[6]_net_1\, 
        \APB3_RDATA_2_i[6]\, \APB3_RDATA_1rs[7]\, 
        \APB3_RDATA_1[7]_net_1\, \APB3_RDATA_2_i[7]_net_1\, 
        \CoreAPB3_0_APBmslave0_PRDATA[0]\, un1_read_reg_en_3_i, 
        \APB3_RDATA_2[0]\, \CoreAPB3_0_APBmslave0_PRDATA[2]\, 
        N_68_i, \CoreAPB3_0_APBmslave0_PRDATA[4]\, 
        \APB3_RDATA_2[4]\, \APB3_RDATA_0_sqmuxa_rs\, 
        \CoreAPB3_0_APBmslave0_PRDATArs[1]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[1]\, APB3_RDATA_0_sqmuxa_i, 
        \APB3_RDATA_2[1]\, \CoreAPB3_0_APBmslave0_PRDATArs[3]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[3]\, N_121_i, 
        \RX_packet_depth[0]_net_1\, \RX_packet_depth_s[0]\, 
        N_416_i, \RX_packet_depth[1]_net_1\, 
        \RX_packet_depth_s[1]\, \RX_packet_depth[2]_net_1\, 
        \RX_packet_depth_s[2]\, \RX_packet_depth[3]_net_1\, 
        \RX_packet_depth_s[3]\, \RX_packet_depth[4]_net_1\, 
        \RX_packet_depth_s[4]\, \RX_packet_depth[5]_net_1\, 
        \RX_packet_depth_s[5]\, \RX_packet_depth[6]_net_1\, 
        \RX_packet_depth_s[6]\, \RX_packet_depth[7]_net_1\, 
        \RX_packet_depth_s[7]_net_1\, RX_packet_depth_s_271_FCO, 
        \RX_packet_depth_cry[0]_net_1\, 
        \RX_packet_depth_cry[1]_net_1\, 
        \RX_packet_depth_cry[2]_net_1\, 
        \RX_packet_depth_cry[3]_net_1\, 
        \RX_packet_depth_cry[4]_net_1\, 
        \RX_packet_depth_cry[5]_net_1\, 
        \RX_packet_depth_cry[6]_net_1\, N_363, 
        \APB3_RDATA_2_8_i_m2_i_m2_0_0_y0[7]\, 
        \APB3_RDATA_2_8_i_m2_i_m2_0_0_co0[7]\, N_500, 
        \APB3_RDATA_2_9_0_0_y0[4]\, \APB3_RDATA_2_9_0_0_co0[4]\, 
        \int_reg[4]\, N_164, \APB3_RDATA_2_7_i_m2_0_0_y0[5]\, 
        \APB3_RDATA_2_7_i_m2_0_0_co0[5]\, N_494, 
        \APB3_RDATA_2_8_0_0_y0[6]\, \APB3_RDATA_2_8_0_0_co0[6]\, 
        N_492, \APB3_RDATA_2_8_0_0_y0[4]\, 
        \APB3_RDATA_2_8_0_0_co0[4]\, N_486, 
        \APB3_RDATA_2_7_0_0_y0[6]\, \APB3_RDATA_2_7_0_0_co0[6]\, 
        N_497, \APB3_RDATA_2_9_0_0_y0[1]\, 
        \APB3_RDATA_2_9_0_0_co0[1]\, \int_reg[1]\, N_489, 
        \APB3_RDATA_2_8_0_0_y0[1]\, \APB3_RDATA_2_8_0_0_co0[1]\, 
        N_161, \APB3_RDATA_2_8_i_m2_0_0_y0[5]\, 
        \APB3_RDATA_2_8_i_m2_0_0_co0[5]\, N_481, 
        \APB3_RDATA_2_7_0_0_y0[1]\, \APB3_RDATA_2_7_0_0_co0[1]\, 
        N_484, \APB3_RDATA_2_7_0_0_y0[4]\, 
        \APB3_RDATA_2_7_0_0_co0[4]\, N_362, 
        \APB3_RDATA_2_7_i_m2_i_m2_0_0_y0[7]\, 
        \APB3_RDATA_2_7_i_m2_i_m2_0_0_co0[7]\, N_162, 
        \APB3_RDATA_2_8_i_m2_0_0_y0[0]\, 
        \APB3_RDATA_2_8_i_m2_0_0_co0[0]\, N_165, 
        \APB3_RDATA_2_7_i_m2_0_0_y0[0]\, 
        \APB3_RDATA_2_7_i_m2_0_0_co0[0]\, N_472, \fifo_MEMRE\, 
        \m14_0_0_1\, N_547, \APB3_RDATA_2_0_i_m2_i_m2_1[7]_net_1\, 
        N_358, m103_1_0, N_104, \APB3_RDATA_2_9_1_1[6]_net_1\, 
        N_502, rx_packet_avail_int, \APB3_RDATA_2_0_1[1]_net_1\, 
        N_423, \APB3_RDATA_2_0_i_m2_1[5]_net_1\, N_177, 
        \APB3_RDATA_2_0_1[6]_net_1\, N_428, 
        \APB3_RDATA_2_0_1[4]_net_1\, N_426, m100_1_0, N_101, 
        \APB3_RDATA_2_0_i_m2_1[0]_net_1\, N_178, 
        \APB3_RDATA_1_RNO_10[3]_net_1\, N_83, 
        \APB3_RDATA_1_RNO_7[2]_net_1\, N_66, 
        \APB3_RDATA_1_RNO_6[3]_net_1\, m47_1_1, 
        \APB3_RDATA_1_RNO_2[3]_net_1\, rx_FIFO_UNDERRUN_int, 
        \APB3_RDATA_1_RNO_8[3]_net_1\, 
        \APB3_RDATA_1_RNO_3[3]_net_1\, 
        \APB3_RDATA_1_RNO_8[2]_net_1\, m59_1_1, 
        \APB3_RDATA_1_RNO_4[2]_net_1\, rx_FIFO_OVERFLOW_int, 
        \APB3_RDATA_1_RNO_10[2]_net_1\, 
        \APB3_RDATA_1_RNO_5[2]_net_1\, \APB3_RDATA_2_am[1]_net_1\, 
        un33_apb3_addr_2, \APB3_RDATA_2_bm[1]_net_1\, 
        \APB3_RDATA_2_am[4]_net_1\, \APB3_RDATA_2_bm[4]_net_1\, 
        N_522, N_512, N_60, N_120, 
        un13_address_low4_reg_en_0_a2_0, un1_apb3_addr_0, \m33_3\, 
        \m33_1\, un1_RX_packet_depthlto7_3, N_299, N_181, N_471, 
        N_71, N_190, N_153, col_detect_int, 
        \APB3_RDATA_2_12_a2_3_0[0]_net_1\, \m33_9\, 
        \APB3_RDATA_2_4_a2_i_0[7]_net_1\, 
        un1_RX_packet_depthlto7_4, \N_480\, \N_6_0\, 
        \un2_apb3_addr_9\, N_329, N_243, N_478, N_540, 
        un1_control_reg_en_2_i_0_0_a2_0_2, un1_apb3_addr_3, 
        \m33_11\, N_26, N_241, N_238, 
        \APB3_RDATA_2_12_1[0]_net_1\, 
        \APB3_RDATA_2_12_0[0]_net_1\, \int_reg[5]\, 
        \APB3_RDATA_2_4_0_1[5]_net_1\, 
        \APB3_RDATA_2_4_0_0[5]_net_1\, \int_reg[7]\, 
        \APB3_RDATA_2_4_0_1[7]_net_1\, 
        \APB3_RDATA_2_4_0_0[7]_net_1\, m33_7, N_559, N_67, N_158, 
        N_159, N_77, N_364, N_388, un10_read_reg_en, 
        \un2_apb3_addr_12\, un25_read_reg_en_0_1, 
        un25_read_reg_en_0_4 : std_logic;

    for all : Interrupts
	Use entity work.Interrupts(DEF_ARCH);
begin 

    consumer_type2_reg(9) <= \consumer_type2_reg[9]\;
    consumer_type2_reg(8) <= \consumer_type2_reg[8]\;
    consumer_type2_reg(7) <= \consumer_type2_reg[7]\;
    consumer_type2_reg(6) <= \consumer_type2_reg[6]\;
    consumer_type2_reg(5) <= \consumer_type2_reg[5]\;
    consumer_type2_reg(4) <= \consumer_type2_reg[4]\;
    consumer_type2_reg(3) <= \consumer_type2_reg[3]\;
    consumer_type2_reg(2) <= \consumer_type2_reg[2]\;
    consumer_type2_reg(1) <= \consumer_type2_reg[1]\;
    consumer_type2_reg(0) <= \consumer_type2_reg[0]\;
    consumer_type3_reg(9) <= \consumer_type3_reg[9]\;
    consumer_type3_reg(8) <= \consumer_type3_reg[8]\;
    consumer_type3_reg(7) <= \consumer_type3_reg[7]\;
    consumer_type3_reg(6) <= \consumer_type3_reg[6]\;
    consumer_type3_reg(5) <= \consumer_type3_reg[5]\;
    consumer_type3_reg(4) <= \consumer_type3_reg[4]\;
    consumer_type3_reg(3) <= \consumer_type3_reg[3]\;
    consumer_type3_reg(2) <= \consumer_type3_reg[2]\;
    consumer_type3_reg(1) <= \consumer_type3_reg[1]\;
    consumer_type3_reg(0) <= \consumer_type3_reg[0]\;
    consumer_type1_reg(9) <= \consumer_type1_reg[9]\;
    consumer_type1_reg(8) <= \consumer_type1_reg[8]\;
    consumer_type1_reg(7) <= \consumer_type1_reg[7]\;
    consumer_type1_reg(6) <= \consumer_type1_reg[6]\;
    consumer_type1_reg(5) <= \consumer_type1_reg[5]\;
    consumer_type1_reg(4) <= \consumer_type1_reg[4]\;
    consumer_type1_reg(3) <= \consumer_type1_reg[3]\;
    consumer_type1_reg(2) <= \consumer_type1_reg[2]\;
    consumer_type1_reg(1) <= \consumer_type1_reg[1]\;
    consumer_type1_reg(0) <= \consumer_type1_reg[0]\;
    consumer_type4_reg(9) <= \consumer_type4_reg[9]\;
    consumer_type4_reg(8) <= \consumer_type4_reg[8]\;
    consumer_type4_reg(7) <= \consumer_type4_reg[7]\;
    consumer_type4_reg(6) <= \consumer_type4_reg[6]\;
    consumer_type4_reg(5) <= \consumer_type4_reg[5]\;
    consumer_type4_reg(4) <= \consumer_type4_reg[4]\;
    consumer_type4_reg(3) <= \consumer_type4_reg[3]\;
    consumer_type4_reg(2) <= \consumer_type4_reg[2]\;
    consumer_type4_reg(1) <= \consumer_type4_reg[1]\;
    consumer_type4_reg(0) <= \consumer_type4_reg[0]\;
    N_6_0 <= \N_6_0\;
    N_480 <= \N_480\;
    fifo_MEMRE <= \fifo_MEMRE\;
    un25_read_reg_en <= \un25_read_reg_en\;
    RX_FIFO_rd_en <= \RX_FIFO_rd_en\;
    TX_FIFO_RST <= \TX_FIFO_RST\;
    start_tx_FIFO <= \start_tx_FIFO\;
    internal_loopback <= \internal_loopback\;
    CoreAPB3_0_APBmslave0_PREADY <= 
        \CoreAPB3_0_APBmslave0_PREADY\;
    un2_apb3_addr_13 <= un2_apb3_addr_13_net_1;
    N_386_i_i <= \N_386_i_i\;

    \control_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_105, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \control_reg[0]_net_1\);
    
    \address_low2_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[2]\);
    
    \WRITE_REGISTER_ENABLE_PROC.un1_apb3_addr_0\ : CFG2
      generic map(INIT => x"2")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => un1_apb3_addr_0);
    
    \APB3_RDATA_1_RNIVKVE[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        \CoreAPB3_0_APBmslave0_PRDATA[2]\, Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(2));
    
    \APB3_RDATA_2_8_i_m2_0_wmux_0[5]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_2_8_i_m2_0_0_y0[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \consumer_type1_reg[5]\, D => \consumer_type2_reg[5]\, 
        FCI => \APB3_RDATA_2_8_i_m2_0_0_co0[5]\, S => OPEN, Y => 
        N_161, FCO => OPEN);
    
    m33_11 : CFG4
      generic map(INIT => x"1000")

      port map(A => rdiff_bus(4), B => rdiff_bus(5), C => \m33_3\, 
        D => \m33_9\, Y => \m33_11\);
    
    \WRITE_REGISTER_ENABLE_PROC.un21_apb3_addr\ : CFG4
      generic map(INIT => x"0040")

      port map(A => N_71, B => N_26, C => 
        CoreAPB3_0_APBmslave0_PADDR(5), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => un21_apb3_addr);
    
    address_low1_reg_en_RNILKOE1 : CFG3
      generic map(INIT => x"20")

      port map(A => \address_low1_reg_en\, B => 
        \address_high1_reg_en\, C => N_472, Y => 
        un13_address_low1_reg_en);
    
    \APB3_RDATA_2_9[6]\ : CFG4
      generic map(INIT => x"EE72")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \APB3_RDATA_2_9_1_1[6]_net_1\, C => rx_FIFO_rst_reg, D
         => CoreAPB3_0_APBmslave0_PADDR(2), Y => N_502);
    
    \APB3_RDATA_2_8_i_m2_0_0_wmux[0]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \consumer_type1_reg[8]\, D => \consumer_type2_reg[8]\, 
        FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_2_8_i_m2_0_0_y0[0]\, FCO => 
        \APB3_RDATA_2_8_i_m2_0_0_co0[0]\);
    
    \WRITE_REGISTER_ENABLE_PROC.address_low4_reg_en_1\ : CFG2
      generic map(INIT => x"2")

      port map(A => \iAPB3_READY[0]_net_1\, B => 
        \CoreAPB3_0_APBmslave0_PREADY\, Y => 
        address_low4_reg_en_1);
    
    \REG_WRITE_PROC.un13_address_low4_reg_en_0_a2_0\ : CFG2
      generic map(INIT => x"4")

      port map(A => \address_high4_reg_en\, B => 
        \address_low4_reg_en\, Y => 
        un13_address_low4_reg_en_0_a2_0);
    
    \RX_PACKET_DEPTH_STATUS_PROC.un1_RX_packet_depthlto7_3\ : 
        CFG2
      generic map(INIT => x"1")

      port map(A => \RX_packet_depth[6]_net_1\, B => 
        \RX_packet_depth[7]_net_1\, Y => 
        un1_RX_packet_depthlto7_3);
    
    \scratch_pad_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[2]_net_1\);
    
    \up_EOP_sync[0]\ : SLE
      port map(D => \up_EOP\, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => long_reset_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \up_EOP_sync[0]_net_1\);
    
    \address_low3_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[2]\);
    
    \WRITE_REGISTER_ENABLE_PROC.un29_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"0008")

      port map(A => N_241, B => un33_apb3_addr_2, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => un29_apb3_addr);
    
    \address_low2_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[6]\);
    
    \APB3_RDATA_2_8_0_wmux_0[4]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_2_8_0_0_y0[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \consumer_type1_reg[4]\, D => \consumer_type2_reg[4]\, 
        FCI => \APB3_RDATA_2_8_0_0_co0[4]\, S => OPEN, Y => N_492, 
        FCO => OPEN);
    
    \APB3_RDATA_1_RNI1NVE[4]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        \CoreAPB3_0_APBmslave0_PRDATA[4]\, Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(4));
    
    \address_low3_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[6]\);
    
    \APB3_RDATA_1_RNO_0[2]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => N_104, C
         => N_66, Y => N_67);
    
    \un2_apb3_addr_13\ : CFG3
      generic map(INIT => x"10")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(1), B => 
        CoreAPB3_0_APBmslave0_PADDR(0), C => \un2_apb3_addr_12\, 
        Y => un2_apb3_addr_13_net_1);
    
    \RX_packet_depth_cry[0]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[0]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        RX_packet_depth_s_271_FCO, S => \RX_packet_depth_s[0]\, Y
         => OPEN, FCO => \RX_packet_depth_cry[0]_net_1\);
    
    read_reg_en_RNIV7T01_0 : CFG1
      generic map(INIT => "01")

      port map(A => N_386_i, Y => \N_386_i_i\);
    
    address_high2_reg_en_RNINGTG : CFG3
      generic map(INIT => x"01")

      port map(A => \address_low1_reg_en\, B => 
        \address_high1_reg_en\, C => \address_high2_reg_en\, Y
         => N_478);
    
    \control_reg_RNO_2[5]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \write_scratch_reg_en\, B => 
        \int_mask_reg_en\, Y => N_471);
    
    \address_low1_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[7]\);
    
    address_low3_reg_en_RNIFRQC2 : CFG3
      generic map(INIT => x"80")

      port map(A => N_559, B => \address_low3_reg_en\, C => N_472, 
        Y => un13_address_low3_reg_en);
    
    address_low2_reg_en_RNI1H422 : CFG3
      generic map(INIT => x"80")

      port map(A => \address_low2_reg_en\, B => N_478, C => N_472, 
        Y => un13_address_low2_reg_en);
    
    \APB3_RDATA_2_11[6]\ : CFG3
      generic map(INIT => x"47")

      port map(A => N_494, B => CoreAPB3_0_APBmslave0_PADDR(5), C
         => N_502, Y => N_522);
    
    \APB3_RDATA_1_RNO[2]\ : CFG3
      generic map(INIT => x"27")

      port map(A => un33_apb3_addr_2, B => N_67, C => N_60, Y => 
        N_68_i);
    
    un2_apb3_addr_9 : CFG3
      generic map(INIT => x"01")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(7), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        CoreAPB3_0_APBmslave0_PADDR(5), Y => \un2_apb3_addr_9\);
    
    \APB3_RDATA_1_RNITIVE[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        \CoreAPB3_0_APBmslave0_PRDATA[0]\, Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(0));
    
    \address_low2_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[4]\);
    
    \APB3_RDATA_2_9_0_0_wmux[4]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => \internal_loopback\, 
        D => \int_reg[4]\, FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_2_9_0_0_y0[4]\, FCO => 
        \APB3_RDATA_2_9_0_0_co0[4]\);
    
    \address_low4_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[4]\);
    
    \APB3_RDATA_2_0_i_m2_1[5]\ : CFG4
      generic map(INIT => x"0F27")

      port map(A => re_pulse_d1, B => RDATA_r(5), C => 
        RDATA_int(5), D => RE_d1, Y => 
        \APB3_RDATA_2_0_i_m2_1[5]_net_1\);
    
    \APB3_RDATA_2_0_i_m2_1[0]\ : CFG4
      generic map(INIT => x"0F27")

      port map(A => re_pulse_d1, B => RDATA_r(0), C => 
        RDATA_int(0), D => RE_d1, Y => 
        \APB3_RDATA_2_0_i_m2_1[0]_net_1\);
    
    \RX_packet_depth_cry[2]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[2]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[1]_net_1\, S => 
        \RX_packet_depth_s[2]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[2]_net_1\);
    
    APB3_RDATA_2_sn_m4_0_a2_0_a2 : CFG2
      generic map(INIT => x"1")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => un33_apb3_addr_2);
    
    \APB3_RDATA_1_RNO_6[2]\ : CFG4
      generic map(INIT => x"0F27")

      port map(A => re_pulse_d1, B => RDATA_r(2), C => 
        RDATA_int(2), D => RE_d1, Y => m103_1_0);
    
    \scratch_pad_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[3]_net_1\);
    
    \APB3_RDATA_2_10_i_m2[5]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => N_177, C
         => N_164, Y => N_158);
    
    \RX_packet_depth[5]\ : SLE
      port map(D => \RX_packet_depth_s[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_416_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[5]_net_1\);
    
    \APB3_RDATA_2_12_a2_3_0[0]\ : CFG3
      generic map(INIT => x"04")

      port map(A => \i_int_mask_reg[0]_net_1\, B => 
        col_detect_int, C => CoreAPB3_0_APBmslave0_PADDR(3), Y
         => \APB3_RDATA_2_12_a2_3_0[0]_net_1\);
    
    \address_high3_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high3_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type3_reg[8]\);
    
    \i_int_mask_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_int_mask_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \i_int_mask_reg[1]_net_1\);
    
    \APB3_RDATA_2_9_0_wmux_0[1]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_2_9_0_0_y0[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \i_int_mask_reg[1]_net_1\, D => RX_FIFO_Full, FCI => 
        \APB3_RDATA_2_9_0_0_co0[1]\, S => OPEN, Y => N_497, FCO
         => OPEN);
    
    \APB3_RDATA_1_RNI71CJ[1]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \APB3_RDATA_0_sqmuxa_rs\, B => 
        \CoreAPB3_0_APBmslave0_PRDATArs[1]\, C => N_386_i_set, Y
         => \CoreAPB3_0_APBmslave0_PRDATA[1]\);
    
    \address_high4_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high4_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high4_reg[2]_net_1\);
    
    \RX_packet_depth[4]\ : SLE
      port map(D => \RX_packet_depth_s[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_416_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[4]_net_1\);
    
    address_high2_reg_en : SLE
      port map(D => address_low4_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un21_apb3_addr, ALn => 
        N_209_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \address_high2_reg_en\);
    
    \WRITE_REGISTER_ENABLE_PROC.un33_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => N_241, B => un33_apb3_addr_2, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => un33_apb3_addr);
    
    \APB3_RDATA_1_RNI4MQI[5]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => N_386_i_rs, B => \APB3_RDATA_1rs[5]\, C => 
        \un2_apb3_addr_13_set\, Y => \APB3_RDATA_1[5]_net_1\);
    
    \APB3_RDATA_2_9_0_0_wmux[1]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => external_loopback, D
         => \int_reg[1]\, FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_2_9_0_0_y0[1]\, FCO => 
        \APB3_RDATA_2_9_0_0_co0[1]\);
    
    \APB3_RDATA_1_RNO_8[2]\ : CFG4
      generic map(INIT => x"F305")

      port map(A => \control_reg[2]_net_1\, B => 
        \i_int_mask_reg[2]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => 
        \APB3_RDATA_1_RNO_8[2]_net_1\);
    
    \REG_READ_PROC.un25_read_reg_en_0_4\ : CFG4
      generic map(INIT => x"FEFC")

      port map(A => N_26, B => un29_apb3_addr, C => 
        un25_read_reg_en_0_1, D => CoreAPB3_0_APBmslave0_PADDR(4), 
        Y => un25_read_reg_en_0_4);
    
    \APB3_RDATA_2_0_i_m2_i_m2_1[7]\ : CFG4
      generic map(INIT => x"0F27")

      port map(A => re_pulse_d1, B => RDATA_r(7), C => 
        RDATA_int(7), D => RE_d1, Y => 
        \APB3_RDATA_2_0_i_m2_i_m2_1[7]_net_1\);
    
    read_reg_en_RNIV7T01 : CFG3
      generic map(INIT => x"3B")

      port map(A => long_reset, B => \read_reg_en\, C => N_540, Y
         => N_386_i);
    
    RX_packet_depth_status_RNO : CFG4
      generic map(INIT => x"EFFF")

      port map(A => \RX_packet_depth[5]_net_1\, B => 
        \RX_packet_depth[4]_net_1\, C => 
        un1_RX_packet_depthlto7_4, D => un1_RX_packet_depthlto7_3, 
        Y => un1_RX_packet_depth_i);
    
    \PROCESSOR_EOP_READ_PROC.un53_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \read_reg_en\, B => 
        \CoreAPB3_0_APBmslave0_PREADY\, C => N_357, D => 
        un45_apb3_addr, Y => un53_apb3_addr);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    RX_packet_depth_s_271 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => rx_packet_complt, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => RX_packet_depth_s_271_FCO);
    
    \address_high2_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high2_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high2_reg[7]_net_1\);
    
    \RX_packet_depth_cry[1]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[1]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[0]_net_1\, S => 
        \RX_packet_depth_s[1]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[1]_net_1\);
    
    \APB3_RDATA_2_7_i_m2_0_0_wmux[0]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \consumer_type3_reg[8]\, D => \consumer_type3_reg[0]\, 
        FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_2_7_i_m2_0_0_y0[0]\, FCO => 
        \APB3_RDATA_2_7_i_m2_0_0_co0[0]\);
    
    \APB3_RDATA_2_12_m2[0]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => RX_FIFO_Empty, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \i_int_mask_reg[0]_net_1\, Y => N_153);
    
    \address_high3_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high3_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high3_reg[5]_net_1\);
    
    \APB3_RDATA_1[6]\ : SLE
      port map(D => \APB3_RDATA_2_i[6]\, CLK => 
        \un25_read_reg_en\, EN => VCC_net_1, ALn => \N_386_i_i\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => VCC_net_1, Q => \APB3_RDATA_1rs[6]\);
    
    \WRITE_REGISTER_ENABLE_PROC.apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => un33_apb3_addr_2, D
         => N_26, Y => apb3_addr);
    
    \m35\ : CFG4
      generic map(INIT => x"D0F0")

      port map(A => iTX_FIFO_rd_en, B => TX_FIFO_Empty, C => 
        REN_d1, D => byte_clk_en, Y => m35);
    
    \APB3_RDATA_1_RNO_5[2]\ : CFG4
      generic map(INIT => x"4C6E")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \APB3_RDATA_1_RNO_10[2]_net_1\, C => 
        \consumer_type2_reg[2]\, D => \consumer_type1_reg[2]\, Y
         => \APB3_RDATA_1_RNO_5[2]_net_1\);
    
    \RX_packet_depth[7]\ : SLE
      port map(D => \RX_packet_depth_s[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_416_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[7]_net_1\);
    
    \APB3_RDATA_2_0_1[6]\ : CFG4
      generic map(INIT => x"0F27")

      port map(A => re_pulse_d1, B => RDATA_r(6), C => 
        RDATA_int(6), D => RE_d1, Y => 
        \APB3_RDATA_2_0_1[6]_net_1\);
    
    \APB3_RDATA_2_i[7]\ : CFG4
      generic map(INIT => x"0105")

      port map(A => \APB3_RDATA_2_4_0_1[7]_net_1\, B => 
        un33_apb3_addr_2, C => \APB3_RDATA_2_4_0_0[7]_net_1\, D
         => N_364, Y => \APB3_RDATA_2_i[7]_net_1\);
    
    iRX_FIFO_rd_en_RNIJFNA : CFG3
      generic map(INIT => x"A6")

      port map(A => REN_d1_0, B => \RX_FIFO_rd_en\, C => 
        RX_FIFO_Empty, Y => N_314_i_i);
    
    \APB3_RDATA_2_8_0_wmux_0[6]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_2_8_0_0_y0[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \consumer_type1_reg[6]\, D => \consumer_type2_reg[6]\, 
        FCI => \APB3_RDATA_2_8_0_0_co0[6]\, S => OPEN, Y => N_494, 
        FCO => OPEN);
    
    \APB3_RDATA_2_8_0_0_wmux[6]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \address_high1_reg[6]_net_1\, D => 
        \address_high2_reg[6]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_2_8_0_0_y0[6]\, FCO => 
        \APB3_RDATA_2_8_0_0_co0[6]\);
    
    m1 : CFG3
      generic map(INIT => x"08")

      port map(A => byte_clk_en, B => iTX_FIFO_rd_en, C => 
        TX_FIFO_Empty, Y => \fifo_MEMRE\);
    
    \RX_packet_depth_cry[5]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[5]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[4]_net_1\, S => 
        \RX_packet_depth_s[5]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[5]_net_1\);
    
    \address_low1_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[1]\);
    
    \control_reg_RNO[5]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(5), B => 
        \control_reg_en\, Y => N_82_i);
    
    \address_high3_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high3_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high3_reg[3]_net_1\);
    
    \address_high4_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high4_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high4_reg[5]_net_1\);
    
    \APB3_RDATA_2_12[0]\ : CFG4
      generic map(INIT => x"FEFC")

      port map(A => un33_apb3_addr_2, B => 
        \APB3_RDATA_2_12_1[0]_net_1\, C => 
        \APB3_RDATA_2_12_0[0]_net_1\, D => N_159, Y => 
        \APB3_RDATA_2[0]\);
    
    \WRITE_REGISTER_ENABLE_PROC.un37_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"0800")

      port map(A => N_241, B => un33_apb3_addr_2, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => un37_apb3_addr);
    
    \APB3_RDATA_2_0_i_m2[5]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \APB3_RDATA_2_0_i_m2_1[5]_net_1\, B => 
        \scratch_pad_reg[5]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_177);
    
    \scratch_pad_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[1]_net_1\);
    
    \i_int_mask_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_int_mask_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \i_int_mask_reg[6]_net_1\);
    
    \iAPB3_READY_RNI02ML[1]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => CoreAPB3_0_APBmslave0_PREADYrs, B => 
        un5_apb3_rst_rs, C => long_reset_set, Y => 
        \CoreAPB3_0_APBmslave0_PREADY\);
    
    \control_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_105, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => rx_FIFO_rst_reg);
    
    \APB3_RDATA_2_ns[4]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_2_am[4]_net_1\, B => 
        un33_apb3_addr_2, C => \APB3_RDATA_2_bm[4]_net_1\, Y => 
        \APB3_RDATA_2[4]\);
    
    \address_high3_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high3_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type3_reg[9]\);
    
    \APB3_RDATA_2_4_0_0[7]\ : CFG4
      generic map(INIT => x"CC50")

      port map(A => \APB3_RDATA_2_4_a2_i_0[7]_net_1\, B => N_363, 
        C => CoreAPB3_0_APBmslave0_PADDR(4), D => 
        CoreAPB3_0_APBmslave0_PADDR(5), Y => 
        \APB3_RDATA_2_4_0_0[7]_net_1\);
    
    \APB3_RDATA_2_7_i_m2_i_m2_0_wmux_0[7]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_2_7_i_m2_i_m2_0_0_y0[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \address_high4_reg[7]_net_1\, D => 
        \consumer_type4_reg[7]\, FCI => 
        \APB3_RDATA_2_7_i_m2_i_m2_0_0_co0[7]\, S => OPEN, Y => 
        N_362, FCO => OPEN);
    
    \APB3_RDATA_2_bm[4]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => N_426, C
         => N_484, Y => \APB3_RDATA_2_bm[4]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un25_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => N_299, B => N_26, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => un25_apb3_addr);
    
    iTX_FIFO_wr_en : SLE
      port map(D => address_low4_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un1_apb3_addr, ALn => 
        N_209_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => TX_FIFO_wr_en);
    
    \APB3_RDATA_2_am[4]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => N_492, C
         => N_500, Y => \APB3_RDATA_2_am[4]_net_1\);
    
    \APB3_RDATA_1_RNIK7VM[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        \CoreAPB3_0_APBmslave0_PRDATA[1]\, Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(1));
    
    \up_EOP_sync[1]\ : SLE
      port map(D => \up_EOP_sync[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \up_EOP_sync[1]_net_1\);
    
    \APB3_RDATA_2_7_0_0_wmux[6]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \address_high3_reg[6]_net_1\, D => 
        \consumer_type3_reg[6]\, FCI => VCC_net_1, S => OPEN, Y
         => \APB3_RDATA_2_7_0_0_y0[6]\, FCO => 
        \APB3_RDATA_2_7_0_0_co0[6]\);
    
    read_reg_en : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => N_384_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \read_reg_en\);
    
    \RX_packet_depth[3]\ : SLE
      port map(D => \RX_packet_depth_s[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_416_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[3]_net_1\);
    
    \address_high3_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high3_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high3_reg[2]_net_1\);
    
    \address_high1_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high1_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high1_reg[6]_net_1\);
    
    \APB3_RDATA_1_RNO_9[2]\ : CFG2
      generic map(INIT => x"2")

      port map(A => rx_FIFO_OVERFLOW_int, B => 
        \i_int_mask_reg[2]_net_1\, Y => m59_1_1);
    
    \APB3_RDATA_1_RNIJUDM[7]\ : CFG2
      generic map(INIT => x"2")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        \APB3_RDATA_1[7]_net_1\, Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(7));
    
    \address_low2_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[1]\);
    
    \WRITE_REGISTER_ENABLE_PROC.un5_apb3_addr_0_a2\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_26, B => N_243, Y => un5_apb3_addr);
    
    \address_low4_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[3]\);
    
    \iAPB3_READY[1]\ : SLE
      port map(D => \iAPB3_READY[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        un5_apb3_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAPB3_0_APBmslave0_PREADYrs);
    
    address_high4_reg_en : SLE
      port map(D => address_low4_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un37_apb3_addr, ALn => 
        N_209_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \address_high4_reg_en\);
    
    \address_low3_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[5]\);
    
    \APB3_RDATA_1_RNO_1[3]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => N_101, C
         => N_83, Y => N_77);
    
    \APB3_RDATA_2_8_0_wmux_0[1]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_2_8_0_0_y0[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \consumer_type1_reg[1]\, D => \consumer_type2_reg[1]\, 
        FCI => \APB3_RDATA_2_8_0_0_co0[1]\, S => OPEN, Y => N_489, 
        FCO => OPEN);
    
    \address_high3_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high3_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high3_reg[4]_net_1\);
    
    \address_high2_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high2_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type2_reg[8]\);
    
    address_high1_reg_en : SLE
      port map(D => address_low4_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_apb3_addr, ALn => 
        N_209_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \address_high1_reg_en\);
    
    \address_low1_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[3]\);
    
    \address_high1_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high1_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high1_reg[5]_net_1\);
    
    \address_high2_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high2_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high2_reg[4]_net_1\);
    
    \APB3_RDATA_1_RNO[3]\ : CFG3
      generic map(INIT => x"1B")

      port map(A => un33_apb3_addr_2, B => N_120, C => N_77, Y
         => N_121_i);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \READY_DELAY_PROC.un5_apb3_rst_rs\ : SLE
      port map(D => VCC_net_1, CLK => long_reset, EN => VCC_net_1, 
        ALn => un5_apb3_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => VCC_net_1, Q => un5_apb3_rst_rs);
    
    \control_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_105, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \control_reg[2]_net_1\);
    
    \APB3_RDATA_2_9_1_1[6]\ : CFG3
      generic map(INIT => x"45")

      port map(A => \i_int_mask_reg[6]_net_1\, B => 
        rx_packet_avail_int, C => CoreAPB3_0_APBmslave0_PADDR(2), 
        Y => \APB3_RDATA_2_9_1_1[6]_net_1\);
    
    \control_reg_RNIS9SH1[1]\ : CFG3
      generic map(INIT => x"02")

      port map(A => DRVR_EN_c, B => tx_packet_complt, C => 
        \N_6_0\, Y => \control_reg_RNIS9SH1[1]_net_1\);
    
    \APB3_RDATA_1_RNO_4[2]\ : CFG4
      generic map(INIT => x"4C6E")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \APB3_RDATA_1_RNO_8[2]_net_1\, C => TX_FIFO_Empty, D => 
        m59_1_1, Y => \APB3_RDATA_1_RNO_4[2]_net_1\);
    
    \i_int_mask_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_int_mask_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \i_int_mask_reg[7]_net_1\);
    
    \address_high4_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high4_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high4_reg[4]_net_1\);
    
    m14_0_0_a5 : CFG3
      generic map(INIT => x"02")

      port map(A => N_190, B => TX_PreAmble, C => un19_tx_dataen, 
        Y => N_547);
    
    \APB3_RDATA_2_8_i_m2_0_wmux_0[0]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_2_8_i_m2_0_0_y0[0]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \consumer_type1_reg[0]\, D => \consumer_type2_reg[0]\, 
        FCI => \APB3_RDATA_2_8_i_m2_0_0_co0[0]\, S => OPEN, Y => 
        N_162, FCO => OPEN);
    
    \address_low4_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[5]\);
    
    \APB3_RDATA_2_7_i_m2_0_wmux_0[0]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_2_7_i_m2_0_0_y0[0]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \consumer_type4_reg[8]\, D => \consumer_type4_reg[0]\, 
        FCI => \APB3_RDATA_2_7_i_m2_0_0_co0[0]\, S => OPEN, Y => 
        N_165, FCO => OPEN);
    
    up_EOP : SLE
      port map(D => un53_apb3_addr, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \up_EOP\);
    
    address_low3_reg_en : SLE
      port map(D => address_low4_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un33_apb3_addr, ALn => 
        N_209_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \address_low3_reg_en\);
    
    \APB3_RDATA_2_i[5]\ : CFG4
      generic map(INIT => x"0105")

      port map(A => \APB3_RDATA_2_4_0_1[5]_net_1\, B => 
        un33_apb3_addr_2, C => \APB3_RDATA_2_4_0_0[5]_net_1\, D
         => N_158, Y => \APB3_RDATA_2_i[5]_net_1\);
    
    \APB3_RDATA_1[2]\ : SLE
      port map(D => N_68_i, CLK => \un25_read_reg_en\, EN => 
        VCC_net_1, ALn => un1_read_reg_en_3_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q
         => \CoreAPB3_0_APBmslave0_PRDATA[2]\);
    
    iRX_FIFO_rd_en_RNIA8LS : CFG4
      generic map(INIT => x"00E0")

      port map(A => rdiff_bus_cry_0_Y_0, B => \RX_FIFO_rd_en\, C
         => \m33_1\, D => rdiff_bus(1), Y => m33_7);
    
    \address_low1_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[0]\);
    
    APB3_RDATA_0_sqmuxa_rs : SLE
      port map(D => VCC_net_1, CLK => N_386_i, EN => VCC_net_1, 
        ALn => APB3_RDATA_0_sqmuxa_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \APB3_RDATA_0_sqmuxa_rs\);
    
    \address_low1_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[2]\);
    
    \RX_packet_depth[6]\ : SLE
      port map(D => \RX_packet_depth_s[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_416_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[6]_net_1\);
    
    \scratch_pad_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[6]_net_1\);
    
    \APB3_RDATA_1[0]\ : SLE
      port map(D => \APB3_RDATA_2[0]\, CLK => \un25_read_reg_en\, 
        EN => VCC_net_1, ALn => un1_read_reg_en_3_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        VCC_net_1, Q => \CoreAPB3_0_APBmslave0_PRDATA[0]\);
    
    \address_high3_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high3_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high3_reg[6]_net_1\);
    
    \REG_READ_PROC.un25_read_reg_en_0_a2_0\ : CFG3
      generic map(INIT => x"02")

      port map(A => N_26, B => CoreAPB3_0_APBmslave0_PADDR(5), C
         => CoreAPB3_0_APBmslave0_PADDR(3), Y => N_388);
    
    \address_low4_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[6]\);
    
    \APB3_RDATA_2_8_i_m2_0_0_wmux[5]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \address_high1_reg[5]_net_1\, D => 
        \address_high2_reg[5]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_2_8_i_m2_0_0_y0[5]\, FCO => 
        \APB3_RDATA_2_8_i_m2_0_0_co0[5]\);
    
    m14_0_0_1 : CFG4
      generic map(INIT => x"2722")

      port map(A => TX_PreAmble, B => tx_preamble_pat_en, C => 
        un19_tx_dataen, D => BIT_CLK, Y => \m14_0_0_1\);
    
    iRX_FIFO_rd_en_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \iAPB3_READY[0]_net_1\, Y => 
        \iAPB3_READY_i[0]\);
    
    \address_low4_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[0]\);
    
    \APB3_RDATA_1_RNO_3[3]\ : CFG4
      generic map(INIT => x"4C6E")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \APB3_RDATA_1_RNO_8[3]_net_1\, C => 
        \consumer_type2_reg[3]\, D => \consumer_type1_reg[3]\, Y
         => \APB3_RDATA_1_RNO_3[3]_net_1\);
    
    \RX_packet_depth[1]\ : SLE
      port map(D => \RX_packet_depth_s[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_416_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[1]_net_1\);
    
    m33_9 : CFG4
      generic map(INIT => x"0001")

      port map(A => rdiff_bus(8), B => rdiff_bus(9), C => 
        rdiff_bus(10), D => rdiff_bus(11), Y => \m33_9\);
    
    \WRITE_REGISTER_ENABLE_PROC.un1_apb3_addr_3\ : CFG4
      generic map(INIT => x"0004")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        un1_apb3_addr_0, C => CoreAPB3_0_APBmslave0_PADDR(4), D
         => CoreAPB3_0_APBmslave0_PADDR(5), Y => un1_apb3_addr_3);
    
    iRX_FIFO_rd_en : SLE
      port map(D => \iAPB3_READY_i[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un45_apb3_addr, ALn => 
        N_384_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \RX_FIFO_rd_en\);
    
    \address_high1_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high1_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type1_reg[9]\);
    
    \address_high2_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high2_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high2_reg[3]_net_1\);
    
    int_mask_reg_en : SLE
      port map(D => address_low4_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un9_apb3_addr, ALn => 
        N_209_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \int_mask_reg_en\);
    
    \address_low1_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[6]\);
    
    \APB3_RDATA_2_0[4]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \APB3_RDATA_2_0_1[4]_net_1\, B => 
        \scratch_pad_reg[4]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_426);
    
    \APB3_RDATA_1_RNIM9VM[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        \CoreAPB3_0_APBmslave0_PRDATA[3]\, Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(3));
    
    \address_low3_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[1]\);
    
    control_reg_en : SLE
      port map(D => address_low4_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un5_apb3_addr, ALn => 
        N_209_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \control_reg_en\);
    
    \APB3_RDATA_1_RNO_5[3]\ : CFG4
      generic map(INIT => x"46CE")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \APB3_RDATA_1_RNO_10[3]_net_1\, C => 
        \address_high4_reg[3]_net_1\, D => 
        \consumer_type4_reg[3]\, Y => N_83);
    
    address_high3_reg_en_RNI4KU71 : CFG3
      generic map(INIT => x"04")

      port map(A => \address_low2_reg_en\, B => N_478, C => 
        \address_high3_reg_en\, Y => N_559);
    
    \REG_WRITE_PROC.un13_address_low4_reg_en_0_a2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => un13_address_low4_reg_en_0_a2_0, B => 
        \address_low3_reg_en\, C => N_559, D => N_472, Y => 
        un13_address_low4_reg_en);
    
    \APB3_RDATA_2_4_a2_i_0[7]\ : CFG3
      generic map(INIT => x"57")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \i_int_mask_reg[7]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => 
        \APB3_RDATA_2_4_a2_i_0[7]_net_1\);
    
    RX_packet_depth_status : SLE
      port map(D => un1_RX_packet_depth_i, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \RX_packet_depth_status\);
    
    \READ_FIFO_ENABLE_PROC.un45_apb3_addr_0_a2_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => un33_apb3_addr_2, D
         => N_26, Y => un45_apb3_addr);
    
    \RX_packet_depth[2]\ : SLE
      port map(D => \RX_packet_depth_s[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_416_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[2]_net_1\);
    
    \scratch_pad_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[7]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un9_apb3_addr_0_a2_0_i\ : CFG3
      generic map(INIT => x"BF")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_329);
    
    \APB3_RDATA_1[1]\ : SLE
      port map(D => \APB3_RDATA_2[1]\, CLK => \un25_read_reg_en\, 
        EN => VCC_net_1, ALn => APB3_RDATA_0_sqmuxa_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        VCC_net_1, Q => \CoreAPB3_0_APBmslave0_PRDATArs[1]\);
    
    \address_low2_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[3]\);
    
    address_high4_reg_en_RNIUB1P2 : CFG4
      generic map(INIT => x"2000")

      port map(A => \address_high4_reg_en\, B => 
        \address_low3_reg_en\, C => N_472, D => N_559, Y => 
        un13_address_high4_reg_en);
    
    \APB3_RDATA_2_4_o2[5]\ : CFG2
      generic map(INIT => x"E")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \i_int_mask_reg[5]_net_1\, Y => N_181);
    
    \APB3_RDATA_2_0_1[1]\ : CFG4
      generic map(INIT => x"0F27")

      port map(A => re_pulse_d1, B => RDATA_r(1), C => 
        RDATA_int(1), D => RE_d1, Y => 
        \APB3_RDATA_2_0_1[1]_net_1\);
    
    \APB3_RDATA_1_RNO_8[3]\ : CFG4
      generic map(INIT => x"F035")

      port map(A => \address_high1_reg[3]_net_1\, B => 
        \address_high2_reg[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => 
        \APB3_RDATA_1_RNO_8[3]_net_1\);
    
    \address_low3_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[0]\);
    
    \address_high1_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high1_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type1_reg[8]\);
    
    \RX_packet_depth[0]\ : SLE
      port map(D => \RX_packet_depth_s[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_416_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[0]_net_1\);
    
    \APB3_RDATA_1[5]\ : SLE
      port map(D => \APB3_RDATA_2_i[5]_net_1\, CLK => 
        \un25_read_reg_en\, EN => VCC_net_1, ALn => \N_386_i_i\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => VCC_net_1, Q => \APB3_RDATA_1rs[5]\);
    
    \address_low4_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[1]\);
    
    \address_high4_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high4_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high4_reg[7]_net_1\);
    
    \APB3_RDATA_1_RNIHSDM[5]\ : CFG2
      generic map(INIT => x"2")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        \APB3_RDATA_1[5]_net_1\, Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(5));
    
    \SYNC2_APB3_CLK_PROC.RX_FIFO_RST_1\ : CFG2
      generic map(INIT => x"E")

      port map(A => RX_EarlyTerm, B => rx_FIFO_rst_reg, Y => 
        RX_FIFO_RST_1);
    
    \REG_READ_PROC.un25_read_reg_en_0\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => un41_apb3_addr, B => un37_apb3_addr, C => 
        un33_apb3_addr, D => un25_read_reg_en_0_4, Y => 
        \un25_read_reg_en\);
    
    \WRITE_REGISTER_ENABLE_PROC.un9_apb3_addr_1_i\ : CFG2
      generic map(INIT => x"7")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_71);
    
    \APB3_RDATA_1_RNO_2[3]\ : CFG4
      generic map(INIT => x"4C6E")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \APB3_RDATA_1_RNO_6[3]_net_1\, C => TX_FIFO_Full, D => 
        m47_1_1, Y => \APB3_RDATA_1_RNO_2[3]_net_1\);
    
    \APB3_RDATA_2_10_i_m2[0]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => N_178, C
         => N_165, Y => N_159);
    
    \APB3_RDATA_2_ns[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_2_am[1]_net_1\, B => 
        un33_apb3_addr_2, C => \APB3_RDATA_2_bm[1]_net_1\, Y => 
        \APB3_RDATA_2[1]\);
    
    m14_0_0_m2_0 : CFG3
      generic map(INIT => x"2E")

      port map(A => p2s_data_0, B => TX_PostAmble_d1, C => 
        BIT_CLK, Y => N_190);
    
    \APB3_RDATA_2_i_ns[6]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un33_apb3_addr_2, B => N_522, C => N_512, Y
         => \APB3_RDATA_2_i[6]\);
    
    \APB3_RDATA_2_7_0_wmux_0[4]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_2_7_0_0_y0[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \address_high4_reg[4]_net_1\, D => 
        \consumer_type4_reg[4]\, FCI => 
        \APB3_RDATA_2_7_0_0_co0[4]\, S => OPEN, Y => N_484, FCO
         => OPEN);
    
    \control_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_105, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => external_loopback);
    
    \address_high2_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high2_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high2_reg[2]_net_1\);
    
    \address_high2_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high2_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high2_reg[6]_net_1\);
    
    \iAPB3_READY[0]\ : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => un5_apb3_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \iAPB3_READYrs[0]\);
    
    \APB3_RDATA_1_RNO_9[3]\ : CFG4
      generic map(INIT => x"0F27")

      port map(A => re_pulse_d1, B => RDATA_r(3), C => 
        RDATA_int(3), D => RE_d1, Y => m100_1_0);
    
    \iRX_FIFO_rd_en_RNIJFNA_0\ : CFG3
      generic map(INIT => x"A2")

      port map(A => REN_d1_0, B => \RX_FIFO_rd_en\, C => 
        RX_FIFO_Empty, Y => iRX_FIFO_rd_en_RNIJFNA_0);
    
    \WRITE_REGISTER_ENABLE_PROC.un41_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => N_241, B => un33_apb3_addr_2, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => un41_apb3_addr);
    
    N_384_i : CFG2
      generic map(INIT => x"2")

      port map(A => N_540, B => long_reset, Y => N_384_i_i);
    
    \APB3_RDATA_2_0_i_m2[0]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \APB3_RDATA_2_0_i_m2_1[0]_net_1\, B => 
        \scratch_pad_reg[0]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_178);
    
    \APB3_RDATA_2_8_i_m2_i_m2_0_0_wmux[7]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \address_high1_reg[7]_net_1\, D => 
        \address_high2_reg[7]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_2_8_i_m2_i_m2_0_0_y0[7]\, FCO => 
        \APB3_RDATA_2_8_i_m2_i_m2_0_0_co0[7]\);
    
    \address_low1_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[4]\);
    
    \i_int_mask_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_int_mask_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \i_int_mask_reg[5]_net_1\);
    
    \address_low4_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[2]\);
    
    m14_0_0 : CFG4
      generic map(INIT => x"FF36")

      port map(A => p2s_data_0, B => BIT_CLK, C => \m14_0_0_1\, D
         => N_547, Y => MANCHESTER_OUT_5);
    
    address_low4_reg_en : SLE
      port map(D => address_low4_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un41_apb3_addr, ALn => 
        N_209_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \address_low4_reg_en\);
    
    m33_1 : CFG2
      generic map(INIT => x"1")

      port map(A => rdiff_bus(2), B => rdiff_bus(3), Y => \m33_1\);
    
    \APB3_RDATA_2_0_i_m2_i_m2[7]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \APB3_RDATA_2_0_i_m2_i_m2_1[7]_net_1\, B => 
        \scratch_pad_reg[7]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_358);
    
    \APB3_RDATA_1_RNO_0[3]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_1_RNO_2[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \APB3_RDATA_1_RNO_3[3]_net_1\, Y => N_120);
    
    un1_read_reg_en_3 : CFG4
      generic map(INIT => x"0C04")

      port map(A => long_reset, B => \read_reg_en\, C => 
        un10_read_reg_en, D => N_540, Y => un1_read_reg_en_3_i);
    
    address_low2_reg_en : SLE
      port map(D => address_low4_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un25_apb3_addr, ALn => 
        N_209_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \address_low2_reg_en\);
    
    \control_reg_RNO_0[5]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => N_559, B => un1_control_reg_en_2_i_0_0_a2_0_2, 
        C => \address_low3_reg_en\, D => control_reg_105, Y => 
        un1_control_reg_en_2_i_0);
    
    \address_low2_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[7]\);
    
    address_high3_reg_en : SLE
      port map(D => address_low4_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un29_apb3_addr, ALn => 
        N_209_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \address_high3_reg_en\);
    
    \APB3_RDATA_2_8_i_m2_i_m2_0_wmux_0[7]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_2_8_i_m2_i_m2_0_0_y0[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \consumer_type1_reg[7]\, D => \consumer_type2_reg[7]\, 
        FCI => \APB3_RDATA_2_8_i_m2_i_m2_0_0_co0[7]\, S => OPEN, 
        Y => N_363, FCO => OPEN);
    
    \APB3_RDATA_2_10_i_m2_i_m2[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_362, B => CoreAPB3_0_APBmslave0_PADDR(6), C
         => N_358, Y => N_364);
    
    \APB3_RDATA_2_0[6]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \APB3_RDATA_2_0_1[6]_net_1\, B => 
        \scratch_pad_reg[6]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_428);
    
    \REG_READ_PROC.un25_read_reg_en_0_1\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_26, B => un33_apb3_addr_2, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => N_388, Y => 
        un25_read_reg_en_0_1);
    
    \N_209_i\ : CFG4
      generic map(INIT => x"0080")

      port map(A => CoreAPB3_0_APBmslave0_PWRITE, B => 
        CoreAPB3_0_APBmslave0_PSELx, C => 
        CoreAPB3_0_APBmslave0_PENABLE, D => long_reset, Y => 
        N_209_i);
    
    \APB3_RDATA_2_10[6]\ : CFG3
      generic map(INIT => x"1B")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => N_428, C
         => N_486, Y => N_512);
    
    \WRITE_REGISTER_ENABLE_PROC.un25_apb3_addr_0_a2_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_299);
    
    \control_reg_RNO_1[5]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => TX_PreAmble, B => \address_low4_reg_en\, C
         => \address_high4_reg_en\, D => N_471, Y => 
        un1_control_reg_en_2_i_0_0_a2_0_2);
    
    \APB3_RDATA_2_bm[1]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => N_423, C
         => N_481, Y => \APB3_RDATA_2_bm[1]_net_1\);
    
    \READY_DELAY_PROC.un5_apb3_rst_0_a2_0_a2\ : CFG3
      generic map(INIT => x"F8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        CoreAPB3_0_APBmslave0_PENABLE, C => long_reset, Y => 
        un5_apb3_rst_i);
    
    \APB3_RDATA_2_am[1]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => N_489, C
         => N_497, Y => \APB3_RDATA_2_am[1]_net_1\);
    
    \RX_packet_depth_cry[6]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[6]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[5]_net_1\, S => 
        \RX_packet_depth_s[6]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[6]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un13_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"0008")

      port map(A => N_299, B => N_26, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => un13_apb3_addr);
    
    \APB3_RDATA_2_12_0[0]\ : CFG4
      generic map(INIT => x"D5C0")

      port map(A => N_329, B => N_162, C => 
        CoreAPB3_0_APBmslave0_PADDR(5), D => N_153, Y => 
        \APB3_RDATA_2_12_0[0]_net_1\);
    
    un2_apb3_addr_12 : CFG4
      generic map(INIT => x"8002")

      port map(A => \un2_apb3_addr_9\, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \un2_apb3_addr_12\);
    
    \address_high4_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high4_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high4_reg[6]_net_1\);
    
    \scratch_pad_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[0]_net_1\);
    
    \APB3_RDATA_1_RNIITDM[6]\ : CFG2
      generic map(INIT => x"2")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        \APB3_RDATA_1[6]_net_1\, Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(6));
    
    \APB3_RDATA_2_7_i_m2_0_wmux_0[5]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_2_7_i_m2_0_0_y0[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \address_high4_reg[5]_net_1\, D => 
        \consumer_type4_reg[5]\, FCI => 
        \APB3_RDATA_2_7_i_m2_0_0_co0[5]\, S => OPEN, Y => N_164, 
        FCO => OPEN);
    
    \i_int_mask_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_int_mask_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \i_int_mask_reg[3]_net_1\);
    
    \address_low1_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[5]\);
    
    \address_high2_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high2_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high2_reg[5]_net_1\);
    
    \REG_WRITE_PROC.un13_address_high1_reg_en_0_a2_0_a2\ : CFG4
      generic map(INIT => x"0004")

      port map(A => \int_mask_reg_en\, B => 
        \address_high1_reg_en\, C => \control_reg_en\, D => 
        \write_scratch_reg_en\, Y => un13_address_high1_reg_en);
    
    address_high3_reg_en_RNIFQLA2 : CFG4
      generic map(INIT => x"4000")

      port map(A => \address_low2_reg_en\, B => 
        \address_high3_reg_en\, C => N_472, D => N_478, Y => 
        un13_address_high3_reg_en);
    
    \address_high3_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high3_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high3_reg[7]_net_1\);
    
    \m34\ : CFG2
      generic map(INIT => x"6")

      port map(A => \fifo_MEMRE\, B => REN_d1, Y => m34);
    
    \up_EOP_sync_RNIOGPQ[2]\ : CFG3
      generic map(INIT => x"9C")

      port map(A => \up_EOP_sync[1]_net_1\, B => rx_packet_complt, 
        C => \up_EOP_sync[2]_net_1\, Y => N_416_i);
    
    \APB3_RDATA_1_RNO_10[2]\ : CFG4
      generic map(INIT => x"F035")

      port map(A => \address_high1_reg[2]_net_1\, B => 
        \address_high2_reg[2]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => 
        \APB3_RDATA_1_RNO_10[2]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un9_apb3_addr_0_a2\ : CFG3
      generic map(INIT => x"04")

      port map(A => N_329, B => N_26, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => un9_apb3_addr);
    
    un2_apb3_addr_13_set : SLE
      port map(D => GND_net_1, CLK => \un25_read_reg_en\, EN => 
        VCC_net_1, ALn => un2_apb3_addr_13_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q
         => \un2_apb3_addr_13_set\);
    
    write_scratch_reg_en : SLE
      port map(D => address_low4_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => apb3_addr, ALn => 
        N_209_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \write_scratch_reg_en\);
    
    \RX_PACKET_DEPTH_STATUS_PROC.un1_RX_packet_depthlto7_4\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \RX_packet_depth[3]_net_1\, B => 
        \RX_packet_depth[2]_net_1\, C => 
        \RX_packet_depth[1]_net_1\, D => 
        \RX_packet_depth[0]_net_1\, Y => 
        un1_RX_packet_depthlto7_4);
    
    INTERRUPT_INST : Interrupts
      port map(CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), 
        CoreAPB3_0_APBmslave0_PADDR(5) => 
        CoreAPB3_0_APBmslave0_PADDR(5), 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        CoreAPB3_0_APBmslave0_PADDR(4), 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(3), 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        CoreAPB3_0_APBmslave0_PADDR(2), i_int_mask_reg(7) => 
        \i_int_mask_reg[7]_net_1\, i_int_mask_reg(6) => 
        \i_int_mask_reg[6]_net_1\, i_int_mask_reg(5) => 
        \i_int_mask_reg[5]_net_1\, i_int_mask_reg(4) => 
        \i_int_mask_reg[4]_net_1\, i_int_mask_reg(3) => 
        \i_int_mask_reg[3]_net_1\, i_int_mask_reg(2) => 
        \i_int_mask_reg[2]_net_1\, i_int_mask_reg(1) => 
        \i_int_mask_reg[1]_net_1\, i_int_mask_reg(0) => 
        \i_int_mask_reg[0]_net_1\, int_reg_6 => \int_reg[7]\, 
        int_reg_3 => \int_reg[4]\, int_reg_0 => \int_reg[1]\, 
        int_reg_4 => \int_reg[5]\, N_26 => N_26, 
        CommsFPGA_top_0_INT => CommsFPGA_top_0_INT, N_238 => 
        N_238, long_reset => long_reset, CommsFPGA_CCC_0_LOCK => 
        CommsFPGA_CCC_0_LOCK, write_reg_en => \write_reg_en\, 
        un29_int_reg_clr => un29_int_reg_clr, N_480_rs => 
        N_480_rs, rx_CRC_error_set => rx_CRC_error_set, 
        un33_int_reg_clr => un33_int_reg_clr, col_detect_int => 
        col_detect_int, N_480_rs_0 => N_480_rs_0, 
        TX_collision_detect_set => TX_collision_detect_set, 
        rx_packet_complt => rx_packet_complt, un9_int_reg_clr => 
        un9_int_reg_clr, rx_packet_avail_int => 
        rx_packet_avail_int, rx_packet_complt_set => 
        rx_packet_complt_set, un13_int_reg_clr => 
        un13_int_reg_clr, N_480_rs_1 => N_480_rs_1, 
        TX_FIFO_UNDERRUN_set => TX_FIFO_UNDERRUN_set, 
        un17_int_reg_clr => un17_int_reg_clr, N_480_rs_2 => 
        N_480_rs_2, TX_FIFO_OVERFLOW_set => TX_FIFO_OVERFLOW_set, 
        un21_int_reg_clr => un21_int_reg_clr, 
        rx_FIFO_UNDERRUN_int => rx_FIFO_UNDERRUN_int, N_480_rs_3
         => N_480_rs_3, RX_FIFO_UNDERRUN_set => 
        RX_FIFO_UNDERRUN_set, un25_int_reg_clr => 
        un25_int_reg_clr, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, rx_FIFO_OVERFLOW_int => 
        rx_FIFO_OVERFLOW_int, N_480_rs_4 => N_480_rs_4, 
        RX_FIFO_OVERFLOW_set => RX_FIFO_OVERFLOW_set, 
        tx_packet_complt => tx_packet_complt, CommsFPGA_CCC_0_GL0
         => CommsFPGA_CCC_0_GL0, N_480_i => N_480_i, N_480 => 
        \N_480\, N_9_0_i_i => N_9_0_i_i);
    
    \control_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_105, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \TX_FIFO_RST\);
    
    \address_high4_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high4_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type4_reg[8]\);
    
    \address_low4_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[7]\);
    
    \i_int_mask_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_int_mask_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \i_int_mask_reg[0]_net_1\);
    
    m36 : CFG2
      generic map(INIT => x"8")

      port map(A => TX_FIFO_rd_en, B => TX_FIFO_Empty, Y => 
        un2_re_p_0);
    
    \scratch_pad_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[4]_net_1\);
    
    int_mask_reg_en_RNIB6N21 : CFG3
      generic map(INIT => x"01")

      port map(A => \write_scratch_reg_en\, B => 
        \int_mask_reg_en\, C => \control_reg_en\, Y => N_472);
    
    \APB3_RDATA_1_RNO_7[2]\ : CFG4
      generic map(INIT => x"F035")

      port map(A => \address_high3_reg[2]_net_1\, B => 
        \address_high4_reg[2]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => 
        \APB3_RDATA_1_RNO_7[2]_net_1\);
    
    \APB3_RDATA_1_RNO_4[3]\ : CFG3
      generic map(INIT => x"A3")

      port map(A => m100_1_0, B => \scratch_pad_reg[3]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), Y => N_101);
    
    \RX_packet_depth_cry[4]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[4]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[3]_net_1\, S => 
        \RX_packet_depth_s[4]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[4]_net_1\);
    
    \APB3_RDATA_1[4]\ : SLE
      port map(D => \APB3_RDATA_2[4]\, CLK => \un25_read_reg_en\, 
        EN => VCC_net_1, ALn => un1_read_reg_en_3_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        VCC_net_1, Q => \CoreAPB3_0_APBmslave0_PRDATA[4]\);
    
    \RX_packet_depth_cry[3]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[3]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[2]_net_1\, S => 
        \RX_packet_depth_s[3]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[3]_net_1\);
    
    \APB3_RDATA_2_0_1[4]\ : CFG4
      generic map(INIT => x"0F27")

      port map(A => re_pulse_d1, B => RDATA_r(4), C => 
        RDATA_int(4), D => RE_d1, Y => 
        \APB3_RDATA_2_0_1[4]_net_1\);
    
    \address_low2_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[0]\);
    
    \APB3_RDATA_2_7_0_wmux_0[6]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_2_7_0_0_y0[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \address_high4_reg[6]_net_1\, D => 
        \consumer_type4_reg[6]\, FCI => 
        \APB3_RDATA_2_7_0_0_co0[6]\, S => OPEN, Y => N_486, FCO
         => OPEN);
    
    \address_low3_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[3]\);
    
    \APB3_RDATA_2_7_i_m2_i_m2_0_0_wmux[7]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \address_high3_reg[7]_net_1\, D => 
        \consumer_type3_reg[7]\, FCI => VCC_net_1, S => OPEN, Y
         => \APB3_RDATA_2_7_i_m2_i_m2_0_0_y0[7]\, FCO => 
        \APB3_RDATA_2_7_i_m2_i_m2_0_0_co0[7]\);
    
    \WRITE_REGISTER_ENABLE_PROC.un17_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => N_299, B => N_26, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => un17_apb3_addr);
    
    \REG_READ_PROC.un10_read_reg_en_0_a2\ : CFG4
      generic map(INIT => x"0008")

      port map(A => N_26, B => un33_apb3_addr_2, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => un10_read_reg_en);
    
    \control_reg_RNIS9SH1_0[1]\ : CLKINT
      port map(A => \control_reg_RNIS9SH1[1]_net_1\, Y => 
        N_106_mux_i_i);
    
    \APB3_RDATA_2_12_1[0]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \APB3_RDATA_2_12_a2_3_0[0]_net_1\, B => 
        \control_reg[0]_net_1\, C => N_243, D => N_238, Y => 
        \APB3_RDATA_2_12_1[0]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un1_apb3_addr\ : CFG4
      generic map(INIT => x"0100")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(7), B => 
        CoreAPB3_0_APBmslave0_PADDR(0), C => 
        CoreAPB3_0_APBmslave0_PADDR(1), D => un1_apb3_addr_3, Y
         => un1_apb3_addr);
    
    iRX_FIFO_rd_en_RNI4O78 : CFG2
      generic map(INIT => x"8")

      port map(A => \RX_FIFO_rd_en\, B => RX_FIFO_Empty, Y => 
        un2_re_p);
    
    \APB3_RDATA_1_RNO_7[3]\ : CFG2
      generic map(INIT => x"2")

      port map(A => rx_FIFO_UNDERRUN_int, B => 
        \i_int_mask_reg[3]_net_1\, Y => m47_1_1);
    
    \address_low3_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[4]\);
    
    \iAPB3_READY_RNIV0ML[0]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \iAPB3_READYrs[0]\, B => un5_apb3_rst_rs, C
         => long_reset_set, Y => \iAPB3_READY[0]_net_1\);
    
    \control_reg[5]\ : SLE
      port map(D => N_82_i, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => un1_control_reg_en_2_i_0, ALn => long_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \start_tx_FIFO\);
    
    \address_low2_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[5]\);
    
    \APB3_RDATA_1[7]\ : SLE
      port map(D => \APB3_RDATA_2_i[7]_net_1\, CLK => 
        \un25_read_reg_en\, EN => VCC_net_1, ALn => \N_386_i_i\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => VCC_net_1, Q => \APB3_RDATA_1rs[7]\);
    
    \address_high4_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high4_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high4_reg[3]_net_1\);
    
    \APB3_RDATA_2_4_0_0[5]\ : CFG4
      generic map(INIT => x"AE0C")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => N_181, C
         => N_329, D => N_161, Y => \APB3_RDATA_2_4_0_0[5]_net_1\);
    
    \APB3_RDATA_1_RNO_3[2]\ : CFG4
      generic map(INIT => x"4C6E")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \APB3_RDATA_1_RNO_7[2]_net_1\, C => 
        \consumer_type4_reg[2]\, D => \consumer_type3_reg[2]\, Y
         => N_66);
    
    \address_high4_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high4_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type4_reg[9]\);
    
    \address_high2_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high2_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \consumer_type2_reg[9]\);
    
    un2_apb3_addr_13_set_RNO : CFG1
      generic map(INIT => "01")

      port map(A => un2_apb3_addr_13_net_1, Y => 
        un2_apb3_addr_13_i);
    
    \APB3_RDATA_2_4_0_1[5]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \int_reg[5]\, B => \start_tx_FIFO\, C => 
        N_243, D => N_238, Y => \APB3_RDATA_2_4_0_1[5]_net_1\);
    
    \APB3_RDATA_1_RNO_10[3]\ : CFG4
      generic map(INIT => x"F035")

      port map(A => \address_high3_reg[3]_net_1\, B => 
        \consumer_type3_reg[3]\, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => 
        \APB3_RDATA_1_RNO_10[3]_net_1\);
    
    apb3_rd_en_i_i_a2 : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PWRITE, B => 
        CoreAPB3_0_APBmslave0_PSELx, C => 
        CoreAPB3_0_APBmslave0_PENABLE, Y => N_540);
    
    address_low1_reg_en : SLE
      port map(D => address_low4_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un17_apb3_addr, ALn => 
        N_209_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \address_low1_reg_en\);
    
    \APB3_RDATA_2_4_0_1[7]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \int_reg[7]\, B => \TX_FIFO_RST\, C => N_243, 
        D => N_238, Y => \APB3_RDATA_2_4_0_1[7]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un5_apb3_addr_0_a2_0\ : CFG4
      generic map(INIT => x"0002")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_243);
    
    \APB3_RDATA_2_7_0_wmux_0[1]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_2_7_0_0_y0[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \consumer_type4_reg[9]\, D => \consumer_type4_reg[1]\, 
        FCI => \APB3_RDATA_2_7_0_0_co0[1]\, S => OPEN, Y => N_481, 
        FCO => OPEN);
    
    \address_low3_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_address_low3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[7]\);
    
    iRX_FIFO_rd_en_RNI4O78_0 : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_rd_en\, B => RX_FIFO_Empty, Y => 
        N_283_i);
    
    \APB3_RDATA_2_0[1]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \APB3_RDATA_2_0_1[1]_net_1\, B => 
        \scratch_pad_reg[1]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_423);
    
    m33_3 : CFG2
      generic map(INIT => x"1")

      port map(A => rdiff_bus(7), B => rdiff_bus(6), Y => \m33_3\);
    
    iRX_FIFO_rd_en_RNI0L4J3 : CFG4
      generic map(INIT => x"1000")

      port map(A => rdiff_bus(12), B => rdiff_bus(13), C => m33_7, 
        D => \m33_11\, Y => empty_r_3);
    
    control_reg_en_RNIVP6K : CFG2
      generic map(INIT => x"4")

      port map(A => \write_scratch_reg_en\, B => \control_reg_en\, 
        Y => control_reg_105);
    
    \APB3_RDATA_2_9_0_wmux_0[4]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_2_9_0_0_y0[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \i_int_mask_reg[4]_net_1\, D => \RX_packet_depth_status\, 
        FCI => \APB3_RDATA_2_9_0_0_co0[4]\, S => OPEN, Y => N_500, 
        FCO => OPEN);
    
    \APB3_RDATA_1_RNO_1[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_1_RNO_4[2]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \APB3_RDATA_1_RNO_5[2]_net_1\, Y => N_60);
    
    \address_high1_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high1_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high1_reg[4]_net_1\);
    
    \APB3_RDATA_2_8_0_0_wmux[4]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \address_high1_reg[4]_net_1\, D => 
        \address_high2_reg[4]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_2_8_0_0_y0[4]\, FCO => 
        \APB3_RDATA_2_8_0_0_co0[4]\);
    
    \APB3_RDATA_2_7_i_m2_0_0_wmux[5]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \address_high3_reg[5]_net_1\, D => 
        \consumer_type3_reg[5]\, FCI => VCC_net_1, S => OPEN, Y
         => \APB3_RDATA_2_7_i_m2_0_0_y0[5]\, FCO => 
        \APB3_RDATA_2_7_i_m2_0_0_co0[5]\);
    
    address_high2_reg_en_RNI2NKJ1 : CFG4
      generic map(INIT => x"0040")

      port map(A => \address_low1_reg_en\, B => 
        \address_high2_reg_en\, C => N_472, D => 
        \address_high1_reg_en\, Y => un13_address_high2_reg_en);
    
    write_reg_en : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => N_209_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \write_reg_en\);
    
    \control_reg_RNIR1VT[1]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \internal_loopback\, B => external_loopback, 
        C => \N_480\, Y => \N_6_0\);
    
    \WRITE_REGISTER_ENABLE_PROC.un21_apb3_addr_2_0_0_a2_0_a2\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(0), B => 
        CoreAPB3_0_APBmslave0_PADDR(1), C => 
        CoreAPB3_0_APBmslave0_PADDR(7), D => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => N_26);
    
    \address_high1_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high1_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high1_reg[3]_net_1\);
    
    \APB3_RDATA_1_RNO_2[2]\ : CFG3
      generic map(INIT => x"A3")

      port map(A => m103_1_0, B => \scratch_pad_reg[2]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), Y => N_104);
    
    \APB3_RDATA_2_8_0_0_wmux[1]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \consumer_type1_reg[9]\, D => \consumer_type2_reg[9]\, 
        FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_2_8_0_0_y0[1]\, FCO => 
        \APB3_RDATA_2_8_0_0_co0[1]\);
    
    \APB3_RDATA_1_RNO_6[3]\ : CFG4
      generic map(INIT => x"F305")

      port map(A => \control_reg[3]_net_1\, B => 
        \i_int_mask_reg[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => 
        \APB3_RDATA_1_RNO_6[3]_net_1\);
    
    \APB3_RDATA_1[3]\ : SLE
      port map(D => N_121_i, CLK => \un25_read_reg_en\, EN => 
        VCC_net_1, ALn => APB3_RDATA_0_sqmuxa_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q
         => \CoreAPB3_0_APBmslave0_PRDATArs[3]\);
    
    \WRITE_REGISTER_ENABLE_PROC.un41_apb3_addr_0_a2_0\ : CFG4
      generic map(INIT => x"0100")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(0), B => 
        CoreAPB3_0_APBmslave0_PADDR(1), C => 
        CoreAPB3_0_APBmslave0_PADDR(7), D => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => N_241);
    
    \i_int_mask_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_int_mask_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \i_int_mask_reg[4]_net_1\);
    
    \REG_WRITE_PROC.un13_int_mask_reg_en_0_a2_0_a2\ : CFG3
      generic map(INIT => x"10")

      port map(A => \control_reg_en\, B => \write_scratch_reg_en\, 
        C => \int_mask_reg_en\, Y => un13_int_mask_reg_en);
    
    \APB3_RDATA_2_7_0_0_wmux[4]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \address_high3_reg[4]_net_1\, D => 
        \consumer_type3_reg[4]\, FCI => VCC_net_1, S => OPEN, Y
         => \APB3_RDATA_2_7_0_0_y0[4]\, FCO => 
        \APB3_RDATA_2_7_0_0_co0[4]\);
    
    \APB3_RDATA_1_RNI6OQI[7]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => N_386_i_rs, B => \APB3_RDATA_1rs[7]\, C => 
        \un2_apb3_addr_13_set\, Y => \APB3_RDATA_1[7]_net_1\);
    
    \APB3_RDATA_1_RNI93CJ[3]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \APB3_RDATA_0_sqmuxa_rs\, B => 
        \CoreAPB3_0_APBmslave0_PRDATArs[3]\, C => N_386_i_set, Y
         => \CoreAPB3_0_APBmslave0_PRDATA[3]\);
    
    \address_high1_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high1_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high1_reg[7]_net_1\);
    
    \RX_packet_depth_s[7]\ : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \RX_packet_depth[7]_net_1\, C
         => rx_packet_complt, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[6]_net_1\, S => 
        \RX_packet_depth_s[7]_net_1\, Y => OPEN, FCO => OPEN);
    
    APB3_RDATA_0_sqmuxa : CFG4
      generic map(INIT => x"3FBF")

      port map(A => long_reset, B => \read_reg_en\, C => 
        un10_read_reg_en, D => N_540, Y => APB3_RDATA_0_sqmuxa_i);
    
    \control_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_105, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \control_reg[3]_net_1\);
    
    \APB3_RDATA_1_RNI5NQI[6]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => N_386_i_rs, B => \APB3_RDATA_1rs[6]\, C => 
        \un2_apb3_addr_13_set\, Y => \APB3_RDATA_1[6]_net_1\);
    
    \i_int_mask_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_int_mask_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \i_int_mask_reg[2]_net_1\);
    
    \scratch_pad_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[5]_net_1\);
    
    \control_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_105, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \internal_loopback\);
    
    \APB3_RDATA_2_7_0_0_wmux[1]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \consumer_type3_reg[9]\, D => \consumer_type3_reg[1]\, 
        FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_2_7_0_0_y0[1]\, FCO => 
        \APB3_RDATA_2_7_0_0_co0[1]\);
    
    \address_high1_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_address_high1_reg_en, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \address_high1_reg[2]_net_1\);
    
    \up_EOP_sync[2]\ : SLE
      port map(D => \up_EOP_sync[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \up_EOP_sync[2]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CommsFPGA_top is

    port( CoreAPB3_0_APBmslave0_PWDATA       : in    std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA_m     : out   std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PADDR        : in    std_logic_vector(7 downto 0);
          DEBOUNCE_IN_c                      : in    std_logic_vector(2 downto 0);
          Y_net_0                            : in    std_logic_vector(3 downto 1);
          DEBOUNCE_OUT_net_0_0               : out   std_logic;
          MANCHESTER_IN_c                    : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY_i_m_i : out   std_logic;
          MANCH_OUT_P_c                      : out   std_logic;
          MANCH_OUT_P_c_i                    : out   std_logic;
          N_209_i_i                          : in    std_logic;
          CoreAPB3_0_APBmslave0_PSELx        : in    std_logic;
          CoreAPB3_0_APBmslave0_PWRITE       : in    std_logic;
          CoreAPB3_0_APBmslave0_PENABLE      : in    std_logic;
          N_209_i                            : out   std_logic;
          DRVR_EN_c                          : out   std_logic;
          CommsFPGA_top_0_INT                : out   std_logic;
          CommsFPGA_CCC_0_LOCK               : in    std_logic;
          DEBOUNCE_OUT_1_c                   : out   std_logic;
          DEBOUNCE_OUT_2_c                   : out   std_logic;
          CommsFPGA_top_0_CAMERA_NODE        : out   std_logic;
          m2s010_som_sb_0_POWER_ON_RESET_N   : in    std_logic;
          m2s010_som_sb_0_GPIO_28_SW_RESET   : in    std_logic;
          CommsFPGA_CCC_0_GL1                : in    std_logic;
          CommsFPGA_CCC_0_GL0                : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz          : in    std_logic
        );

end CommsFPGA_top;

architecture DEF_ARCH of CommsFPGA_top is 

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component TriDebounce
    port( DEBOUNCE_IN_c        : in    std_logic_vector(2 downto 0) := (others => 'U');
          DEBOUNCE_OUT_net_0_0 : out   std_logic;
          DEBOUNCE_OUT_2_c     : out   std_logic;
          DEBOUNCE_OUT_1_c     : out   std_logic;
          BIT_CLK              : in    std_logic := 'U';
          N_480_set            : in    std_logic := 'U';
          N_480                : in    std_logic := 'U'
        );
  end component;

  component ManchesEncoder
    port( manches_in_dly        : in    std_logic_vector(1 downto 0) := (others => 'U');
          RX_FIFO_DIN           : in    std_logic_vector(7 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe_0    : in    std_logic := 'U';
          p2s_data_0            : out   std_logic;
          N_9_0_i_i             : in    std_logic := 'U';
          start_tx_FIFO         : in    std_logic := 'U';
          iTX_FIFO_rd_en        : out   std_logic;
          tx_packet_complt      : out   std_logic;
          TX_PreAmble           : out   std_logic;
          TX_FIFO_Empty         : in    std_logic := 'U';
          TX_FIFO_rd_en         : out   std_logic;
          N_268_i               : out   std_logic;
          TX_collision_detect   : out   std_logic;
          TX_collision_detect_i : out   std_logic;
          N_106_mux_i_i         : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0   : in    std_logic := 'U';
          N_366_i               : in    std_logic := 'U';
          tx_col_detect_en      : out   std_logic;
          N_6_0                 : in    std_logic := 'U';
          DRVR_EN_c             : out   std_logic;
          rx_crc_HighByte_en    : in    std_logic := 'U';
          un19_tx_dataen        : out   std_logic;
          N_517                 : in    std_logic := 'U';
          N_522                 : in    std_logic := 'U';
          N_519                 : in    std_logic := 'U';
          N_518                 : in    std_logic := 'U';
          N_521                 : in    std_logic := 'U';
          N_520                 : in    std_logic := 'U';
          N_228                 : in    std_logic := 'U';
          N_516                 : in    std_logic := 'U';
          tx_preamble_pat_en    : out   std_logic;
          TX_PostAmble_d1       : out   std_logic;
          MANCHESTER_OUT_5      : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL1   : in    std_logic := 'U';
          byte_clk_en           : in    std_logic := 'U';
          BIT_CLK               : in    std_logic := 'U';
          N_480_i               : in    std_logic := 'U';
          MANCH_OUT_P_c_i       : out   std_logic;
          MANCH_OUT_P_c         : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component ManchesDecoder
    port( RX_FIFO_DIN_pipe                   : out   std_logic_vector(8 downto 0);
          consumer_type1_reg                 : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type2_reg                 : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type3_reg                 : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type4_reg                 : in    std_logic_vector(9 downto 0) := (others => 'U');
          RX_FIFO_DIN                        : out   std_logic_vector(7 downto 0);
          manches_in_dly                     : out   std_logic_vector(1 downto 0);
          rx_CRC_error                       : out   std_logic;
          rx_CRC_error_i                     : out   std_logic;
          rx_packet_complt                   : out   std_logic;
          rx_packet_complt_i                 : out   std_logic;
          rx_crc_HighByte_en                 : out   std_logic;
          iRX_FIFO_wr_en                     : out   std_logic;
          RX_InProcess_d1                    : out   std_logic;
          TX_collision_detect                : in    std_logic := 'U';
          tx_col_detect_en                   : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PSELx        : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY       : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY_i_m_i : out   std_logic;
          N_366_i                            : out   std_logic;
          DRVR_EN_c                          : in    std_logic := 'U';
          CommsFPGA_CCC_0_LOCK               : in    std_logic := 'U';
          long_reset                         : in    std_logic := 'U';
          N_480                              : in    std_logic := 'U';
          RX_EarlyTerm                       : out   std_logic;
          CommsFPGA_CCC_0_GL0                : in    std_logic := 'U';
          N_480_i                            : in    std_logic := 'U';
          sampler_clk1x_en                   : out   std_logic;
          MANCH_OUT_P_c                      : in    std_logic := 'U';
          MANCHESTER_IN_c                    : in    std_logic := 'U';
          internal_loopback                  : in    std_logic := 'U';
          N_268_i                            : in    std_logic := 'U'
        );
  end component;

  component FIFOs
    port( RX_FIFO_DIN_pipe             : in    std_logic_vector(8 downto 0) := (others => 'U');
          rdiff_bus                    : out   std_logic_vector(13 downto 1);
          RDATA_int                    : out   std_logic_vector(7 downto 0);
          RDATA_r                      : out   std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          RX_FIFO_UNDERRUN             : out   std_logic;
          RX_FIFO_UNDERRUN_i           : out   std_logic;
          RX_FIFO_OVERFLOW             : out   std_logic;
          RX_FIFO_OVERFLOW_i           : out   std_logic;
          CommsFPGA_CCC_0_GL0          : in    std_logic := 'U';
          RX_FIFO_Empty                : out   std_logic;
          empty_r_3                    : in    std_logic := 'U';
          RX_FIFO_Full                 : out   std_logic;
          un2_re_p_0                   : in    std_logic := 'U';
          rdiff_bus_cry_0_Y_0          : out   std_logic;
          iRX_FIFO_wr_en               : in    std_logic := 'U';
          sampler_clk1x_en             : in    std_logic := 'U';
          RX_InProcess_d1              : in    std_logic := 'U';
          tx_col_detect_en             : in    std_logic := 'U';
          N_357                        : out   std_logic;
          re_pulse_d1                  : out   std_logic;
          RX_FIFO_rd_en                : in    std_logic := 'U';
          RE_d1                        : out   std_logic;
          N_283_i                      : in    std_logic := 'U';
          N_314_i_i                    : in    std_logic := 'U';
          REN_d1_0                     : out   std_logic;
          iRX_FIFO_rd_en_RNIJFNA_0     : in    std_logic := 'U';
          TX_FIFO_UNDERRUN             : out   std_logic;
          TX_FIFO_UNDERRUN_i           : out   std_logic;
          TX_FIFO_OVERFLOW             : out   std_logic;
          TX_FIFO_OVERFLOW_i           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic := 'U';
          un2_re_p                     : in    std_logic := 'U';
          TX_FIFO_Empty                : out   std_logic;
          TX_FIFO_Full                 : out   std_logic;
          TX_FIFO_wr_en                : in    std_logic := 'U';
          N_516                        : out   std_logic;
          N_517                        : out   std_logic;
          N_518                        : out   std_logic;
          N_519                        : out   std_logic;
          N_520                        : out   std_logic;
          N_521                        : out   std_logic;
          N_228                        : out   std_logic;
          N_522                        : out   std_logic;
          TX_FIFO_rd_en                : in    std_logic := 'U';
          fifo_MEMRE                   : in    std_logic := 'U';
          m34                          : in    std_logic := 'U';
          REN_d1                       : out   std_logic;
          m35                          : in    std_logic := 'U';
          BIT_CLK                      : in    std_logic := 'U';
          RX_FIFO_RST                  : in    std_logic := 'U';
          TX_FIFO_RST                  : in    std_logic := 'U';
          N_480                        : in    std_logic := 'U'
        );
  end component;

  component uP_if
    port( rdiff_bus                      : in    std_logic_vector(13 downto 1) := (others => 'U');
          CoreAPB3_0_APBmslave0_PADDR    : in    std_logic_vector(7 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PRDATA_m : out   std_logic_vector(7 downto 0);
          RDATA_int                      : in    std_logic_vector(7 downto 0) := (others => 'U');
          RDATA_r                        : in    std_logic_vector(7 downto 0) := (others => 'U');
          consumer_type2_reg             : out   std_logic_vector(9 downto 0);
          consumer_type3_reg             : out   std_logic_vector(9 downto 0);
          consumer_type1_reg             : out   std_logic_vector(9 downto 0);
          consumer_type4_reg             : out   std_logic_vector(9 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA   : in    std_logic_vector(7 downto 0) := (others => 'U');
          p2s_data_0                     : in    std_logic := 'U';
          N_9_0_i_i                      : out   std_logic;
          N_480_i                        : out   std_logic;
          RX_FIFO_OVERFLOW_set           : in    std_logic := 'U';
          N_480_rs_4                     : in    std_logic := 'U';
          un25_int_reg_clr               : out   std_logic;
          RX_FIFO_UNDERRUN_set           : in    std_logic := 'U';
          N_480_rs_3                     : in    std_logic := 'U';
          un21_int_reg_clr               : out   std_logic;
          TX_FIFO_OVERFLOW_set           : in    std_logic := 'U';
          N_480_rs_2                     : in    std_logic := 'U';
          un17_int_reg_clr               : out   std_logic;
          TX_FIFO_UNDERRUN_set           : in    std_logic := 'U';
          N_480_rs_1                     : in    std_logic := 'U';
          un13_int_reg_clr               : out   std_logic;
          rx_packet_complt_set           : in    std_logic := 'U';
          un9_int_reg_clr                : out   std_logic;
          TX_collision_detect_set        : in    std_logic := 'U';
          N_480_rs_0                     : in    std_logic := 'U';
          un33_int_reg_clr               : out   std_logic;
          rx_CRC_error_set               : in    std_logic := 'U';
          N_480_rs                       : in    std_logic := 'U';
          un29_int_reg_clr               : out   std_logic;
          CommsFPGA_CCC_0_LOCK           : in    std_logic := 'U';
          CommsFPGA_top_0_INT            : out   std_logic;
          empty_r_3                      : out   std_logic;
          N_357                          : in    std_logic := 'U';
          tx_packet_complt               : in    std_logic := 'U';
          DRVR_EN_c                      : in    std_logic := 'U';
          N_209_i                        : out   std_logic;
          rdiff_bus_cry_0_Y_0            : in    std_logic := 'U';
          N_314_i_i                      : out   std_logic;
          m34                            : out   std_logic;
          un2_re_p_0                     : out   std_logic;
          TX_FIFO_rd_en                  : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PENABLE  : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PWRITE   : in    std_logic := 'U';
          iRX_FIFO_rd_en_RNIJFNA_0       : out   std_logic;
          REN_d1_0                       : in    std_logic := 'U';
          N_283_i                        : out   std_logic;
          N_6_0                          : out   std_logic;
          N_480                          : out   std_logic;
          TX_PostAmble_d1                : in    std_logic := 'U';
          RX_FIFO_RST_1                  : out   std_logic;
          RX_EarlyTerm                   : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PSELx    : in    std_logic := 'U';
          un2_re_p                       : out   std_logic;
          RX_FIFO_Empty                  : in    std_logic := 'U';
          TX_FIFO_Full                   : in    std_logic := 'U';
          RE_d1                          : in    std_logic := 'U';
          re_pulse_d1                    : in    std_logic := 'U';
          un19_tx_dataen                 : in    std_logic := 'U';
          tx_preamble_pat_en             : in    std_logic := 'U';
          TX_PreAmble                    : in    std_logic := 'U';
          MANCHESTER_OUT_5               : out   std_logic;
          BIT_CLK                        : in    std_logic := 'U';
          fifo_MEMRE                     : out   std_logic;
          m35                            : out   std_logic;
          byte_clk_en                    : in    std_logic := 'U';
          REN_d1                         : in    std_logic := 'U';
          TX_FIFO_Empty                  : in    std_logic := 'U';
          iTX_FIFO_rd_en                 : in    std_logic := 'U';
          RX_FIFO_Full                   : in    std_logic := 'U';
          rx_packet_complt               : in    std_logic := 'U';
          N_386_i_set                    : in    std_logic := 'U';
          un25_read_reg_en               : out   std_logic;
          N_386_i_rs                     : in    std_logic := 'U';
          TX_FIFO_wr_en                  : out   std_logic;
          N_209_i_i                      : in    std_logic := 'U';
          RX_FIFO_rd_en                  : out   std_logic;
          TX_FIFO_RST                    : out   std_logic;
          start_tx_FIFO                  : out   std_logic;
          internal_loopback              : out   std_logic;
          long_reset                     : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY   : out   std_logic;
          long_reset_set                 : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz      : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0            : in    std_logic := 'U';
          long_reset_i                   : in    std_logic := 'U';
          un2_apb3_addr_13               : out   std_logic;
          N_386_i_i                      : out   std_logic;
          N_106_mux_i_i                  : out   std_logic
        );
  end component;

    signal bd_reset_i, \bd_reset\, \long_reset\, long_reset_0, 
        \BIT_CLK\, BIT_CLK_0, \ClkDivider[0]_net_1\, 
        \ClkDivider_i[0]\, BIT_CLK_i_i, long_reset_i, \N_480_set\, 
        GND_net_1, N_480_i, VCC_net_1, \long_reset_set\, 
        \RX_FIFO_OVERFLOW_set\, RX_FIFO_OVERFLOW_i, 
        un25_int_reg_clr, \N_480_rs_4\, RX_FIFO_OVERFLOW, 
        \RX_FIFO_UNDERRUN_set\, RX_FIFO_UNDERRUN_i, 
        un21_int_reg_clr, \N_480_rs_3\, RX_FIFO_UNDERRUN, 
        \TX_FIFO_OVERFLOW_set\, TX_FIFO_OVERFLOW_i, 
        un17_int_reg_clr, \N_480_rs_2\, TX_FIFO_OVERFLOW, 
        \TX_FIFO_UNDERRUN_set\, TX_FIFO_UNDERRUN_i, 
        un13_int_reg_clr, \N_480_rs_1\, TX_FIFO_UNDERRUN, 
        \rx_packet_complt_set\, rx_packet_complt_i, 
        un9_int_reg_clr, \TX_collision_detect_set\, 
        TX_collision_detect_i, un33_int_reg_clr, \N_480_rs_0\, 
        TX_collision_detect, \rx_CRC_error_set\, rx_CRC_error_i, 
        un29_int_reg_clr, \N_480_rs\, rx_CRC_error, 
        \ClkDivider[1]_net_1\, \ClkDivider_RNO[1]_net_1\, 
        \ClkDivider[2]_net_1\, \ClkDivider_RNO[2]_net_1\, 
        \long_reset_cntr[0]_net_1\, \long_reset_cntr_3[0]_net_1\, 
        \long_reset_cntr[1]_net_1\, \long_reset_cntr_3[1]_net_1\, 
        \long_reset_cntr[2]_net_1\, \long_reset_cntr_3[2]_net_1\, 
        \long_reset_cntr[3]_net_1\, \long_reset_cntr_3[3]_net_1\, 
        \long_reset_cntr[4]_net_1\, \long_reset_cntr_3[4]_net_1\, 
        \long_reset_cntr[5]_net_1\, \long_reset_cntr_3[5]_net_1\, 
        \long_reset_cntr[6]_net_1\, un4_long_reset_cntr_cry_6_S, 
        \long_reset_cntr[7]_net_1\, un4_long_reset_cntr_s_7_S, 
        un2_long_reset_cntr_i, \RX_FIFO_RST\, RX_FIFO_RST_1, 
        \byte_clk_en\, byte_clk_en_1, \N_386_i_rs\, N_386_i_i, 
        un2_apb3_addr_13, \N_386_i_set\, un25_read_reg_en, 
        un4_long_reset_cntr_s_1_277_FCO, 
        \un4_long_reset_cntr_cry_1\, un4_long_reset_cntr_cry_1_S, 
        \un4_long_reset_cntr_cry_2\, un4_long_reset_cntr_cry_2_S, 
        \un4_long_reset_cntr_cry_3\, un4_long_reset_cntr_cry_3_S, 
        \un4_long_reset_cntr_cry_4\, un4_long_reset_cntr_cry_4_S, 
        \un4_long_reset_cntr_cry_5\, un4_long_reset_cntr_cry_5_S, 
        \un4_long_reset_cntr_cry_6\, un2_long_reset_cntr_5, 
        un2_long_reset_cntr_4, N_480, \rdiff_bus[1]\, 
        \rdiff_bus[2]\, \rdiff_bus[3]\, \rdiff_bus[4]\, 
        \rdiff_bus[5]\, \rdiff_bus[6]\, \rdiff_bus[7]\, 
        \rdiff_bus[8]\, \rdiff_bus[9]\, \rdiff_bus[10]\, 
        \rdiff_bus[11]\, \rdiff_bus[12]\, \rdiff_bus[13]\, 
        \RDATA_int[0]\, \RDATA_int[1]\, \RDATA_int[2]\, 
        \RDATA_int[3]\, \RDATA_int[4]\, \RDATA_int[5]\, 
        \RDATA_int[6]\, \RDATA_int[7]\, \RDATA_r[0]\, 
        \RDATA_r[1]\, \RDATA_r[2]\, \RDATA_r[3]\, \RDATA_r[4]\, 
        \RDATA_r[5]\, \RDATA_r[6]\, \RDATA_r[7]\, \p2s_data[7]\, 
        \consumer_type2_reg[0]\, \consumer_type2_reg[1]\, 
        \consumer_type2_reg[2]\, \consumer_type2_reg[3]\, 
        \consumer_type2_reg[4]\, \consumer_type2_reg[5]\, 
        \consumer_type2_reg[6]\, \consumer_type2_reg[7]\, 
        \consumer_type2_reg[8]\, \consumer_type2_reg[9]\, 
        \consumer_type3_reg[0]\, \consumer_type3_reg[1]\, 
        \consumer_type3_reg[2]\, \consumer_type3_reg[3]\, 
        \consumer_type3_reg[4]\, \consumer_type3_reg[5]\, 
        \consumer_type3_reg[6]\, \consumer_type3_reg[7]\, 
        \consumer_type3_reg[8]\, \consumer_type3_reg[9]\, 
        \consumer_type1_reg[0]\, \consumer_type1_reg[1]\, 
        \consumer_type1_reg[2]\, \consumer_type1_reg[3]\, 
        \consumer_type1_reg[4]\, \consumer_type1_reg[5]\, 
        \consumer_type1_reg[6]\, \consumer_type1_reg[7]\, 
        \consumer_type1_reg[8]\, \consumer_type1_reg[9]\, 
        \consumer_type4_reg[0]\, \consumer_type4_reg[1]\, 
        \consumer_type4_reg[2]\, \consumer_type4_reg[3]\, 
        \consumer_type4_reg[4]\, \consumer_type4_reg[5]\, 
        \consumer_type4_reg[6]\, \consumer_type4_reg[7]\, 
        \consumer_type4_reg[8]\, \consumer_type4_reg[9]\, 
        N_9_0_i_i, empty_r_3, N_357, tx_packet_complt, 
        \DRVR_EN_c\, rdiff_bus_cry_0_Y_0, N_314_i_i, m34, 
        un2_re_p, TX_FIFO_rd_en, iRX_FIFO_rd_en_RNIJFNA_0, REN_d1, 
        N_283_i, N_6_0, TX_PostAmble_d1, RX_EarlyTerm, un2_re_p_0, 
        RX_FIFO_Empty, TX_FIFO_Full, RE_d1, re_pulse_d1, 
        un19_tx_dataen, tx_preamble_pat_en, TX_PreAmble, 
        MANCHESTER_OUT_5, fifo_MEMRE, m35, REN_d1_0, 
        TX_FIFO_Empty, iTX_FIFO_rd_en, RX_FIFO_Full, 
        rx_packet_complt, TX_FIFO_wr_en, RX_FIFO_rd_en, 
        TX_FIFO_RST, start_tx_FIFO, internal_loopback, 
        CoreAPB3_0_APBmslave0_PREADY, N_106_mux_i_i, 
        \RX_FIFO_DIN_pipe[0]\, \RX_FIFO_DIN_pipe[1]\, 
        \RX_FIFO_DIN_pipe[2]\, \RX_FIFO_DIN_pipe[3]\, 
        \RX_FIFO_DIN_pipe[4]\, \RX_FIFO_DIN_pipe[5]\, 
        \RX_FIFO_DIN_pipe[6]\, \RX_FIFO_DIN_pipe[7]\, 
        \RX_FIFO_DIN_pipe[8]\, iRX_FIFO_wr_en, sampler_clk1x_en, 
        RX_InProcess_d1, tx_col_detect_en, N_516, N_517, N_518, 
        N_519, N_520, N_521, N_228, N_522, \manches_in_dly[0]\, 
        \manches_in_dly[1]\, \RX_FIFO_DIN[0]\, \RX_FIFO_DIN[1]\, 
        \RX_FIFO_DIN[2]\, \RX_FIFO_DIN[3]\, \RX_FIFO_DIN[4]\, 
        \RX_FIFO_DIN[5]\, \RX_FIFO_DIN[6]\, \RX_FIFO_DIN[7]\, 
        N_268_i, N_366_i, rx_crc_HighByte_en, \MANCH_OUT_P_c\
         : std_logic;

    for all : TriDebounce
	Use entity work.TriDebounce(DEF_ARCH);
    for all : ManchesEncoder
	Use entity work.ManchesEncoder(DEF_ARCH);
    for all : ManchesDecoder
	Use entity work.ManchesDecoder(DEF_ARCH);
    for all : FIFOs
	Use entity work.FIFOs(DEF_ARCH);
    for all : uP_if
	Use entity work.uP_if(DEF_ARCH);
begin 

    MANCH_OUT_P_c <= \MANCH_OUT_P_c\;
    DRVR_EN_c <= \DRVR_EN_c\;

    BIT_CLK_inferred_clock_RNIT9E2 : CLKINT
      port map(A => BIT_CLK_0, Y => \BIT_CLK\);
    
    \long_reset_cntr_3[3]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => un2_long_reset_cntr_4, B => 
        un2_long_reset_cntr_5, C => un4_long_reset_cntr_cry_3_S, 
        Y => \long_reset_cntr_3[3]_net_1\);
    
    bd_reset : CFG2
      generic map(INIT => x"4")

      port map(A => m2s010_som_sb_0_GPIO_28_SW_RESET, B => 
        m2s010_som_sb_0_POWER_ON_RESET_N, Y => \bd_reset\);
    
    \long_reset_cntr[3]\ : SLE
      port map(D => \long_reset_cntr_3[3]_net_1\, CLK => 
        \BIT_CLK\, EN => VCC_net_1, ALn => bd_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[3]_net_1\);
    
    \RESET_DELAY_PROC.un2_long_reset_cntr_4\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \long_reset_cntr[4]_net_1\, B => 
        \long_reset_cntr[3]_net_1\, C => 
        \long_reset_cntr[2]_net_1\, D => 
        \long_reset_cntr[1]_net_1\, Y => un2_long_reset_cntr_4);
    
    \long_reset_cntr[6]\ : SLE
      port map(D => un4_long_reset_cntr_cry_6_S, CLK => \BIT_CLK\, 
        EN => VCC_net_1, ALn => bd_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \long_reset_cntr[6]_net_1\);
    
    \ClkDivider_RNO[2]\ : CFG3
      generic map(INIT => x"6A")

      port map(A => \ClkDivider[2]_net_1\, B => 
        \ClkDivider[1]_net_1\, C => \ClkDivider[0]_net_1\, Y => 
        \ClkDivider_RNO[2]_net_1\);
    
    byte_clk_en : SLE
      port map(D => byte_clk_en_1, CLK => \BIT_CLK\, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \byte_clk_en\);
    
    N_480_rs_2 : SLE
      port map(D => VCC_net_1, CLK => TX_FIFO_OVERFLOW, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \N_480_rs_2\);
    
    long_reset_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => long_reset_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \long_reset_set\);
    
    \ClkDivider_RNO[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \ClkDivider[0]_net_1\, B => 
        \ClkDivider[1]_net_1\, Y => \ClkDivider_RNO[1]_net_1\);
    
    \RESET_DELAY_PROC.un2_long_reset_cntr_5\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \long_reset_cntr[7]_net_1\, B => 
        \long_reset_cntr[6]_net_1\, C => 
        \long_reset_cntr[5]_net_1\, D => 
        \long_reset_cntr[0]_net_1\, Y => un2_long_reset_cntr_5);
    
    N_480_rs_3 : SLE
      port map(D => VCC_net_1, CLK => RX_FIFO_UNDERRUN, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \N_480_rs_3\);
    
    un4_long_reset_cntr_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[2]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_1\, S => 
        un4_long_reset_cntr_cry_2_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_2\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \ID_RES_DECODE_PROC.un4_id_res\ : CFG3
      generic map(INIT => x"08")

      port map(A => Y_net_0(3), B => Y_net_0(2), C => Y_net_0(1), 
        Y => CommsFPGA_top_0_CAMERA_NODE);
    
    N_480_rs_4 : SLE
      port map(D => VCC_net_1, CLK => RX_FIFO_OVERFLOW, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \N_480_rs_4\);
    
    \ClkDivider_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \ClkDivider[0]_net_1\, Y => \ClkDivider_i[0]\);
    
    \long_reset_cntr[5]\ : SLE
      port map(D => \long_reset_cntr_3[5]_net_1\, CLK => 
        \BIT_CLK\, EN => VCC_net_1, ALn => bd_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[5]_net_1\);
    
    rx_packet_complt_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un9_int_reg_clr, ALn => rx_packet_complt_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_packet_complt_set\);
    
    N_386_i_set : SLE
      port map(D => GND_net_1, CLK => un25_read_reg_en, EN => 
        VCC_net_1, ALn => N_386_i_i, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \N_386_i_set\);
    
    TRIPLE_DEBOUNCE_INST : TriDebounce
      port map(DEBOUNCE_IN_c(2) => DEBOUNCE_IN_c(2), 
        DEBOUNCE_IN_c(1) => DEBOUNCE_IN_c(1), DEBOUNCE_IN_c(0)
         => DEBOUNCE_IN_c(0), DEBOUNCE_OUT_net_0_0 => 
        DEBOUNCE_OUT_net_0_0, DEBOUNCE_OUT_2_c => 
        DEBOUNCE_OUT_2_c, DEBOUNCE_OUT_1_c => DEBOUNCE_OUT_1_c, 
        BIT_CLK => \BIT_CLK\, N_480_set => \N_480_set\, N_480 => 
        N_480);
    
    un4_long_reset_cntr_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[3]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_2\, S => 
        un4_long_reset_cntr_cry_3_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_3\);
    
    MANCHESTER_ENCODER_INST : ManchesEncoder
      port map(manches_in_dly(1) => \manches_in_dly[1]\, 
        manches_in_dly(0) => \manches_in_dly[0]\, RX_FIFO_DIN(7)
         => \RX_FIFO_DIN[7]\, RX_FIFO_DIN(6) => \RX_FIFO_DIN[6]\, 
        RX_FIFO_DIN(5) => \RX_FIFO_DIN[5]\, RX_FIFO_DIN(4) => 
        \RX_FIFO_DIN[4]\, RX_FIFO_DIN(3) => \RX_FIFO_DIN[3]\, 
        RX_FIFO_DIN(2) => \RX_FIFO_DIN[2]\, RX_FIFO_DIN(1) => 
        \RX_FIFO_DIN[1]\, RX_FIFO_DIN(0) => \RX_FIFO_DIN[0]\, 
        RX_FIFO_DIN_pipe_0 => \RX_FIFO_DIN_pipe[8]\, p2s_data_0
         => \p2s_data[7]\, N_9_0_i_i => N_9_0_i_i, start_tx_FIFO
         => start_tx_FIFO, iTX_FIFO_rd_en => iTX_FIFO_rd_en, 
        tx_packet_complt => tx_packet_complt, TX_PreAmble => 
        TX_PreAmble, TX_FIFO_Empty => TX_FIFO_Empty, 
        TX_FIFO_rd_en => TX_FIFO_rd_en, N_268_i => N_268_i, 
        TX_collision_detect => TX_collision_detect, 
        TX_collision_detect_i => TX_collision_detect_i, 
        N_106_mux_i_i => N_106_mux_i_i, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, N_366_i => N_366_i, tx_col_detect_en
         => tx_col_detect_en, N_6_0 => N_6_0, DRVR_EN_c => 
        \DRVR_EN_c\, rx_crc_HighByte_en => rx_crc_HighByte_en, 
        un19_tx_dataen => un19_tx_dataen, N_517 => N_517, N_522
         => N_522, N_519 => N_519, N_518 => N_518, N_521 => N_521, 
        N_520 => N_520, N_228 => N_228, N_516 => N_516, 
        tx_preamble_pat_en => tx_preamble_pat_en, TX_PostAmble_d1
         => TX_PostAmble_d1, MANCHESTER_OUT_5 => MANCHESTER_OUT_5, 
        CommsFPGA_CCC_0_GL1 => CommsFPGA_CCC_0_GL1, byte_clk_en
         => \byte_clk_en\, BIT_CLK => \BIT_CLK\, N_480_i => 
        N_480_i, MANCH_OUT_P_c_i => MANCH_OUT_P_c_i, 
        MANCH_OUT_P_c => \MANCH_OUT_P_c\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \SAMPLE_5MHZ_EN_PROC.byte_clk_en_1\ : CFG3
      generic map(INIT => x"08")

      port map(A => \ClkDivider[2]_net_1\, B => 
        \ClkDivider[1]_net_1\, C => \ClkDivider[0]_net_1\, Y => 
        byte_clk_en_1);
    
    \long_reset_cntr[7]\ : SLE
      port map(D => un4_long_reset_cntr_s_7_S, CLK => \BIT_CLK\, 
        EN => VCC_net_1, ALn => bd_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \long_reset_cntr[7]_net_1\);
    
    long_reset : SLE
      port map(D => un2_long_reset_cntr_i, CLK => \BIT_CLK\, EN
         => VCC_net_1, ALn => bd_reset_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        long_reset_0);
    
    TX_FIFO_OVERFLOW_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un17_int_reg_clr, ALn => TX_FIFO_OVERFLOW_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \TX_FIFO_OVERFLOW_set\);
    
    RX_FIFO_OVERFLOW_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un25_int_reg_clr, ALn => RX_FIFO_OVERFLOW_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_OVERFLOW_set\);
    
    un4_long_reset_cntr_s_1_277 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[0]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un4_long_reset_cntr_s_1_277_FCO);
    
    un4_long_reset_cntr_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[4]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_3\, S => 
        un4_long_reset_cntr_cry_4_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_4\);
    
    long_reset_RNO : CFG2
      generic map(INIT => x"7")

      port map(A => un2_long_reset_cntr_5, B => 
        un2_long_reset_cntr_4, Y => un2_long_reset_cntr_i);
    
    BIT_CLK : SLE
      port map(D => BIT_CLK_i_i, CLK => CommsFPGA_CCC_0_GL1, EN
         => VCC_net_1, ALn => bd_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        BIT_CLK_0);
    
    MANCHESTER_DECODER_INST : ManchesDecoder
      port map(RX_FIFO_DIN_pipe(8) => \RX_FIFO_DIN_pipe[8]\, 
        RX_FIFO_DIN_pipe(7) => \RX_FIFO_DIN_pipe[7]\, 
        RX_FIFO_DIN_pipe(6) => \RX_FIFO_DIN_pipe[6]\, 
        RX_FIFO_DIN_pipe(5) => \RX_FIFO_DIN_pipe[5]\, 
        RX_FIFO_DIN_pipe(4) => \RX_FIFO_DIN_pipe[4]\, 
        RX_FIFO_DIN_pipe(3) => \RX_FIFO_DIN_pipe[3]\, 
        RX_FIFO_DIN_pipe(2) => \RX_FIFO_DIN_pipe[2]\, 
        RX_FIFO_DIN_pipe(1) => \RX_FIFO_DIN_pipe[1]\, 
        RX_FIFO_DIN_pipe(0) => \RX_FIFO_DIN_pipe[0]\, 
        consumer_type1_reg(9) => \consumer_type1_reg[9]\, 
        consumer_type1_reg(8) => \consumer_type1_reg[8]\, 
        consumer_type1_reg(7) => \consumer_type1_reg[7]\, 
        consumer_type1_reg(6) => \consumer_type1_reg[6]\, 
        consumer_type1_reg(5) => \consumer_type1_reg[5]\, 
        consumer_type1_reg(4) => \consumer_type1_reg[4]\, 
        consumer_type1_reg(3) => \consumer_type1_reg[3]\, 
        consumer_type1_reg(2) => \consumer_type1_reg[2]\, 
        consumer_type1_reg(1) => \consumer_type1_reg[1]\, 
        consumer_type1_reg(0) => \consumer_type1_reg[0]\, 
        consumer_type2_reg(9) => \consumer_type2_reg[9]\, 
        consumer_type2_reg(8) => \consumer_type2_reg[8]\, 
        consumer_type2_reg(7) => \consumer_type2_reg[7]\, 
        consumer_type2_reg(6) => \consumer_type2_reg[6]\, 
        consumer_type2_reg(5) => \consumer_type2_reg[5]\, 
        consumer_type2_reg(4) => \consumer_type2_reg[4]\, 
        consumer_type2_reg(3) => \consumer_type2_reg[3]\, 
        consumer_type2_reg(2) => \consumer_type2_reg[2]\, 
        consumer_type2_reg(1) => \consumer_type2_reg[1]\, 
        consumer_type2_reg(0) => \consumer_type2_reg[0]\, 
        consumer_type3_reg(9) => \consumer_type3_reg[9]\, 
        consumer_type3_reg(8) => \consumer_type3_reg[8]\, 
        consumer_type3_reg(7) => \consumer_type3_reg[7]\, 
        consumer_type3_reg(6) => \consumer_type3_reg[6]\, 
        consumer_type3_reg(5) => \consumer_type3_reg[5]\, 
        consumer_type3_reg(4) => \consumer_type3_reg[4]\, 
        consumer_type3_reg(3) => \consumer_type3_reg[3]\, 
        consumer_type3_reg(2) => \consumer_type3_reg[2]\, 
        consumer_type3_reg(1) => \consumer_type3_reg[1]\, 
        consumer_type3_reg(0) => \consumer_type3_reg[0]\, 
        consumer_type4_reg(9) => \consumer_type4_reg[9]\, 
        consumer_type4_reg(8) => \consumer_type4_reg[8]\, 
        consumer_type4_reg(7) => \consumer_type4_reg[7]\, 
        consumer_type4_reg(6) => \consumer_type4_reg[6]\, 
        consumer_type4_reg(5) => \consumer_type4_reg[5]\, 
        consumer_type4_reg(4) => \consumer_type4_reg[4]\, 
        consumer_type4_reg(3) => \consumer_type4_reg[3]\, 
        consumer_type4_reg(2) => \consumer_type4_reg[2]\, 
        consumer_type4_reg(1) => \consumer_type4_reg[1]\, 
        consumer_type4_reg(0) => \consumer_type4_reg[0]\, 
        RX_FIFO_DIN(7) => \RX_FIFO_DIN[7]\, RX_FIFO_DIN(6) => 
        \RX_FIFO_DIN[6]\, RX_FIFO_DIN(5) => \RX_FIFO_DIN[5]\, 
        RX_FIFO_DIN(4) => \RX_FIFO_DIN[4]\, RX_FIFO_DIN(3) => 
        \RX_FIFO_DIN[3]\, RX_FIFO_DIN(2) => \RX_FIFO_DIN[2]\, 
        RX_FIFO_DIN(1) => \RX_FIFO_DIN[1]\, RX_FIFO_DIN(0) => 
        \RX_FIFO_DIN[0]\, manches_in_dly(1) => 
        \manches_in_dly[1]\, manches_in_dly(0) => 
        \manches_in_dly[0]\, rx_CRC_error => rx_CRC_error, 
        rx_CRC_error_i => rx_CRC_error_i, rx_packet_complt => 
        rx_packet_complt, rx_packet_complt_i => 
        rx_packet_complt_i, rx_crc_HighByte_en => 
        rx_crc_HighByte_en, iRX_FIFO_wr_en => iRX_FIFO_wr_en, 
        RX_InProcess_d1 => RX_InProcess_d1, TX_collision_detect
         => TX_collision_detect, tx_col_detect_en => 
        tx_col_detect_en, CoreAPB3_0_APBmslave0_PSELx => 
        CoreAPB3_0_APBmslave0_PSELx, CoreAPB3_0_APBmslave0_PREADY
         => CoreAPB3_0_APBmslave0_PREADY, 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, N_366_i => N_366_i, 
        DRVR_EN_c => \DRVR_EN_c\, CommsFPGA_CCC_0_LOCK => 
        CommsFPGA_CCC_0_LOCK, long_reset => \long_reset\, N_480
         => N_480, RX_EarlyTerm => RX_EarlyTerm, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, N_480_i => 
        N_480_i, sampler_clk1x_en => sampler_clk1x_en, 
        MANCH_OUT_P_c => \MANCH_OUT_P_c\, MANCHESTER_IN_c => 
        MANCHESTER_IN_c, internal_loopback => internal_loopback, 
        N_268_i => N_268_i);
    
    \long_reset_cntr_3[2]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => un2_long_reset_cntr_4, B => 
        un2_long_reset_cntr_5, C => un4_long_reset_cntr_cry_2_S, 
        Y => \long_reset_cntr_3[2]_net_1\);
    
    N_480_rs_0 : SLE
      port map(D => VCC_net_1, CLK => TX_collision_detect, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \N_480_rs_0\);
    
    N_480_rs : SLE
      port map(D => VCC_net_1, CLK => rx_CRC_error, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \N_480_rs\);
    
    \long_reset_cntr_3[1]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => un2_long_reset_cntr_4, B => 
        un2_long_reset_cntr_5, C => un4_long_reset_cntr_cry_1_S, 
        Y => \long_reset_cntr_3[1]_net_1\);
    
    un4_long_reset_cntr_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[5]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_4\, S => 
        un4_long_reset_cntr_cry_5_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_5\);
    
    un4_long_reset_cntr_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[6]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_5\, S => 
        un4_long_reset_cntr_cry_6_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_6\);
    
    rx_CRC_error_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un29_int_reg_clr, ALn => rx_CRC_error_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_CRC_error_set\);
    
    BIT_CLK_RNO : CFG1
      generic map(INIT => "01")

      port map(A => BIT_CLK_0, Y => BIT_CLK_i_i);
    
    un4_long_reset_cntr_s_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[7]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_6\, S => 
        un4_long_reset_cntr_s_7_S, Y => OPEN, FCO => OPEN);
    
    long_reset_RNIUA27 : CLKINT
      port map(A => long_reset_0, Y => \long_reset\);
    
    N_480_set : SLE
      port map(D => GND_net_1, CLK => \BIT_CLK\, EN => VCC_net_1, 
        ALn => N_480_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \N_480_set\);
    
    \ClkDivider[2]\ : SLE
      port map(D => \ClkDivider_RNO[2]_net_1\, CLK => \BIT_CLK\, 
        EN => VCC_net_1, ALn => bd_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ClkDivider[2]_net_1\);
    
    un4_long_reset_cntr_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[1]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        un4_long_reset_cntr_s_1_277_FCO, S => 
        un4_long_reset_cntr_cry_1_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_1\);
    
    \long_reset_cntr_3[5]\ : CFG3
      generic map(INIT => x"70")

      port map(A => un2_long_reset_cntr_4, B => 
        un2_long_reset_cntr_5, C => un4_long_reset_cntr_cry_5_S, 
        Y => \long_reset_cntr_3[5]_net_1\);
    
    RX_FIFO_RST : SLE
      port map(D => RX_FIFO_RST_1, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => bd_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_RST\);
    
    \ClkDivider[0]\ : SLE
      port map(D => \ClkDivider_i[0]\, CLK => \BIT_CLK\, EN => 
        VCC_net_1, ALn => bd_reset_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ClkDivider[0]_net_1\);
    
    N_480_rs_1 : SLE
      port map(D => VCC_net_1, CLK => TX_FIFO_UNDERRUN, EN => 
        VCC_net_1, ALn => N_480_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \N_480_rs_1\);
    
    long_reset_RNIUA27_0 : CFG1
      generic map(INIT => "01")

      port map(A => \long_reset\, Y => long_reset_i);
    
    \long_reset_cntr[2]\ : SLE
      port map(D => \long_reset_cntr_3[2]_net_1\, CLK => 
        \BIT_CLK\, EN => VCC_net_1, ALn => bd_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[2]_net_1\);
    
    \long_reset_cntr[1]\ : SLE
      port map(D => \long_reset_cntr_3[1]_net_1\, CLK => 
        \BIT_CLK\, EN => VCC_net_1, ALn => bd_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[1]_net_1\);
    
    \long_reset_cntr_3[0]\ : CFG3
      generic map(INIT => x"B3")

      port map(A => un2_long_reset_cntr_5, B => 
        \long_reset_cntr[0]_net_1\, C => un2_long_reset_cntr_4, Y
         => \long_reset_cntr_3[0]_net_1\);
    
    \long_reset_cntr[0]\ : SLE
      port map(D => \long_reset_cntr_3[0]_net_1\, CLK => 
        \BIT_CLK\, EN => VCC_net_1, ALn => bd_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[0]_net_1\);
    
    TX_FIFO_UNDERRUN_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un13_int_reg_clr, ALn => TX_FIFO_UNDERRUN_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \TX_FIFO_UNDERRUN_set\);
    
    \long_reset_cntr_3[4]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => un2_long_reset_cntr_4, B => 
        un2_long_reset_cntr_5, C => un4_long_reset_cntr_cry_4_S, 
        Y => \long_reset_cntr_3[4]_net_1\);
    
    FIFOS_INST : FIFOs
      port map(RX_FIFO_DIN_pipe(8) => \RX_FIFO_DIN_pipe[8]\, 
        RX_FIFO_DIN_pipe(7) => \RX_FIFO_DIN_pipe[7]\, 
        RX_FIFO_DIN_pipe(6) => \RX_FIFO_DIN_pipe[6]\, 
        RX_FIFO_DIN_pipe(5) => \RX_FIFO_DIN_pipe[5]\, 
        RX_FIFO_DIN_pipe(4) => \RX_FIFO_DIN_pipe[4]\, 
        RX_FIFO_DIN_pipe(3) => \RX_FIFO_DIN_pipe[3]\, 
        RX_FIFO_DIN_pipe(2) => \RX_FIFO_DIN_pipe[2]\, 
        RX_FIFO_DIN_pipe(1) => \RX_FIFO_DIN_pipe[1]\, 
        RX_FIFO_DIN_pipe(0) => \RX_FIFO_DIN_pipe[0]\, 
        rdiff_bus(13) => \rdiff_bus[13]\, rdiff_bus(12) => 
        \rdiff_bus[12]\, rdiff_bus(11) => \rdiff_bus[11]\, 
        rdiff_bus(10) => \rdiff_bus[10]\, rdiff_bus(9) => 
        \rdiff_bus[9]\, rdiff_bus(8) => \rdiff_bus[8]\, 
        rdiff_bus(7) => \rdiff_bus[7]\, rdiff_bus(6) => 
        \rdiff_bus[6]\, rdiff_bus(5) => \rdiff_bus[5]\, 
        rdiff_bus(4) => \rdiff_bus[4]\, rdiff_bus(3) => 
        \rdiff_bus[3]\, rdiff_bus(2) => \rdiff_bus[2]\, 
        rdiff_bus(1) => \rdiff_bus[1]\, RDATA_int(7) => 
        \RDATA_int[7]\, RDATA_int(6) => \RDATA_int[6]\, 
        RDATA_int(5) => \RDATA_int[5]\, RDATA_int(4) => 
        \RDATA_int[4]\, RDATA_int(3) => \RDATA_int[3]\, 
        RDATA_int(2) => \RDATA_int[2]\, RDATA_int(1) => 
        \RDATA_int[1]\, RDATA_int(0) => \RDATA_int[0]\, 
        RDATA_r(7) => \RDATA_r[7]\, RDATA_r(6) => \RDATA_r[6]\, 
        RDATA_r(5) => \RDATA_r[5]\, RDATA_r(4) => \RDATA_r[4]\, 
        RDATA_r(3) => \RDATA_r[3]\, RDATA_r(2) => \RDATA_r[2]\, 
        RDATA_r(1) => \RDATA_r[1]\, RDATA_r(0) => \RDATA_r[0]\, 
        CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), RX_FIFO_UNDERRUN => 
        RX_FIFO_UNDERRUN, RX_FIFO_UNDERRUN_i => 
        RX_FIFO_UNDERRUN_i, RX_FIFO_OVERFLOW => RX_FIFO_OVERFLOW, 
        RX_FIFO_OVERFLOW_i => RX_FIFO_OVERFLOW_i, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, RX_FIFO_Empty
         => RX_FIFO_Empty, empty_r_3 => empty_r_3, RX_FIFO_Full
         => RX_FIFO_Full, un2_re_p_0 => un2_re_p_0, 
        rdiff_bus_cry_0_Y_0 => rdiff_bus_cry_0_Y_0, 
        iRX_FIFO_wr_en => iRX_FIFO_wr_en, sampler_clk1x_en => 
        sampler_clk1x_en, RX_InProcess_d1 => RX_InProcess_d1, 
        tx_col_detect_en => tx_col_detect_en, N_357 => N_357, 
        re_pulse_d1 => re_pulse_d1, RX_FIFO_rd_en => 
        RX_FIFO_rd_en, RE_d1 => RE_d1, N_283_i => N_283_i, 
        N_314_i_i => N_314_i_i, REN_d1_0 => REN_d1, 
        iRX_FIFO_rd_en_RNIJFNA_0 => iRX_FIFO_rd_en_RNIJFNA_0, 
        TX_FIFO_UNDERRUN => TX_FIFO_UNDERRUN, TX_FIFO_UNDERRUN_i
         => TX_FIFO_UNDERRUN_i, TX_FIFO_OVERFLOW => 
        TX_FIFO_OVERFLOW, TX_FIFO_OVERFLOW_i => 
        TX_FIFO_OVERFLOW_i, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, un2_re_p => un2_re_p, 
        TX_FIFO_Empty => TX_FIFO_Empty, TX_FIFO_Full => 
        TX_FIFO_Full, TX_FIFO_wr_en => TX_FIFO_wr_en, N_516 => 
        N_516, N_517 => N_517, N_518 => N_518, N_519 => N_519, 
        N_520 => N_520, N_521 => N_521, N_228 => N_228, N_522 => 
        N_522, TX_FIFO_rd_en => TX_FIFO_rd_en, fifo_MEMRE => 
        fifo_MEMRE, m34 => m34, REN_d1 => REN_d1_0, m35 => m35, 
        BIT_CLK => \BIT_CLK\, RX_FIFO_RST => \RX_FIFO_RST\, 
        TX_FIFO_RST => TX_FIFO_RST, N_480 => N_480);
    
    PROCESSOR_INTERFACE_INST : uP_if
      port map(rdiff_bus(13) => \rdiff_bus[13]\, rdiff_bus(12)
         => \rdiff_bus[12]\, rdiff_bus(11) => \rdiff_bus[11]\, 
        rdiff_bus(10) => \rdiff_bus[10]\, rdiff_bus(9) => 
        \rdiff_bus[9]\, rdiff_bus(8) => \rdiff_bus[8]\, 
        rdiff_bus(7) => \rdiff_bus[7]\, rdiff_bus(6) => 
        \rdiff_bus[6]\, rdiff_bus(5) => \rdiff_bus[5]\, 
        rdiff_bus(4) => \rdiff_bus[4]\, rdiff_bus(3) => 
        \rdiff_bus[3]\, rdiff_bus(2) => \rdiff_bus[2]\, 
        rdiff_bus(1) => \rdiff_bus[1]\, 
        CoreAPB3_0_APBmslave0_PADDR(7) => 
        CoreAPB3_0_APBmslave0_PADDR(7), 
        CoreAPB3_0_APBmslave0_PADDR(6) => 
        CoreAPB3_0_APBmslave0_PADDR(6), 
        CoreAPB3_0_APBmslave0_PADDR(5) => 
        CoreAPB3_0_APBmslave0_PADDR(5), 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        CoreAPB3_0_APBmslave0_PADDR(4), 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(3), 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        CoreAPB3_0_APBmslave0_PADDR(2), 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        CoreAPB3_0_APBmslave0_PADDR(1), 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        CoreAPB3_0_APBmslave0_PADDR(0), 
        CoreAPB3_0_APBmslave0_PRDATA_m(7) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(7), 
        CoreAPB3_0_APBmslave0_PRDATA_m(6) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(6), 
        CoreAPB3_0_APBmslave0_PRDATA_m(5) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(5), 
        CoreAPB3_0_APBmslave0_PRDATA_m(4) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(4), 
        CoreAPB3_0_APBmslave0_PRDATA_m(3) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(3), 
        CoreAPB3_0_APBmslave0_PRDATA_m(2) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(2), 
        CoreAPB3_0_APBmslave0_PRDATA_m(1) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(1), 
        CoreAPB3_0_APBmslave0_PRDATA_m(0) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(0), RDATA_int(7) => 
        \RDATA_int[7]\, RDATA_int(6) => \RDATA_int[6]\, 
        RDATA_int(5) => \RDATA_int[5]\, RDATA_int(4) => 
        \RDATA_int[4]\, RDATA_int(3) => \RDATA_int[3]\, 
        RDATA_int(2) => \RDATA_int[2]\, RDATA_int(1) => 
        \RDATA_int[1]\, RDATA_int(0) => \RDATA_int[0]\, 
        RDATA_r(7) => \RDATA_r[7]\, RDATA_r(6) => \RDATA_r[6]\, 
        RDATA_r(5) => \RDATA_r[5]\, RDATA_r(4) => \RDATA_r[4]\, 
        RDATA_r(3) => \RDATA_r[3]\, RDATA_r(2) => \RDATA_r[2]\, 
        RDATA_r(1) => \RDATA_r[1]\, RDATA_r(0) => \RDATA_r[0]\, 
        consumer_type2_reg(9) => \consumer_type2_reg[9]\, 
        consumer_type2_reg(8) => \consumer_type2_reg[8]\, 
        consumer_type2_reg(7) => \consumer_type2_reg[7]\, 
        consumer_type2_reg(6) => \consumer_type2_reg[6]\, 
        consumer_type2_reg(5) => \consumer_type2_reg[5]\, 
        consumer_type2_reg(4) => \consumer_type2_reg[4]\, 
        consumer_type2_reg(3) => \consumer_type2_reg[3]\, 
        consumer_type2_reg(2) => \consumer_type2_reg[2]\, 
        consumer_type2_reg(1) => \consumer_type2_reg[1]\, 
        consumer_type2_reg(0) => \consumer_type2_reg[0]\, 
        consumer_type3_reg(9) => \consumer_type3_reg[9]\, 
        consumer_type3_reg(8) => \consumer_type3_reg[8]\, 
        consumer_type3_reg(7) => \consumer_type3_reg[7]\, 
        consumer_type3_reg(6) => \consumer_type3_reg[6]\, 
        consumer_type3_reg(5) => \consumer_type3_reg[5]\, 
        consumer_type3_reg(4) => \consumer_type3_reg[4]\, 
        consumer_type3_reg(3) => \consumer_type3_reg[3]\, 
        consumer_type3_reg(2) => \consumer_type3_reg[2]\, 
        consumer_type3_reg(1) => \consumer_type3_reg[1]\, 
        consumer_type3_reg(0) => \consumer_type3_reg[0]\, 
        consumer_type1_reg(9) => \consumer_type1_reg[9]\, 
        consumer_type1_reg(8) => \consumer_type1_reg[8]\, 
        consumer_type1_reg(7) => \consumer_type1_reg[7]\, 
        consumer_type1_reg(6) => \consumer_type1_reg[6]\, 
        consumer_type1_reg(5) => \consumer_type1_reg[5]\, 
        consumer_type1_reg(4) => \consumer_type1_reg[4]\, 
        consumer_type1_reg(3) => \consumer_type1_reg[3]\, 
        consumer_type1_reg(2) => \consumer_type1_reg[2]\, 
        consumer_type1_reg(1) => \consumer_type1_reg[1]\, 
        consumer_type1_reg(0) => \consumer_type1_reg[0]\, 
        consumer_type4_reg(9) => \consumer_type4_reg[9]\, 
        consumer_type4_reg(8) => \consumer_type4_reg[8]\, 
        consumer_type4_reg(7) => \consumer_type4_reg[7]\, 
        consumer_type4_reg(6) => \consumer_type4_reg[6]\, 
        consumer_type4_reg(5) => \consumer_type4_reg[5]\, 
        consumer_type4_reg(4) => \consumer_type4_reg[4]\, 
        consumer_type4_reg(3) => \consumer_type4_reg[3]\, 
        consumer_type4_reg(2) => \consumer_type4_reg[2]\, 
        consumer_type4_reg(1) => \consumer_type4_reg[1]\, 
        consumer_type4_reg(0) => \consumer_type4_reg[0]\, 
        CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), p2s_data_0 => 
        \p2s_data[7]\, N_9_0_i_i => N_9_0_i_i, N_480_i => N_480_i, 
        RX_FIFO_OVERFLOW_set => \RX_FIFO_OVERFLOW_set\, 
        N_480_rs_4 => \N_480_rs_4\, un25_int_reg_clr => 
        un25_int_reg_clr, RX_FIFO_UNDERRUN_set => 
        \RX_FIFO_UNDERRUN_set\, N_480_rs_3 => \N_480_rs_3\, 
        un21_int_reg_clr => un21_int_reg_clr, 
        TX_FIFO_OVERFLOW_set => \TX_FIFO_OVERFLOW_set\, 
        N_480_rs_2 => \N_480_rs_2\, un17_int_reg_clr => 
        un17_int_reg_clr, TX_FIFO_UNDERRUN_set => 
        \TX_FIFO_UNDERRUN_set\, N_480_rs_1 => \N_480_rs_1\, 
        un13_int_reg_clr => un13_int_reg_clr, 
        rx_packet_complt_set => \rx_packet_complt_set\, 
        un9_int_reg_clr => un9_int_reg_clr, 
        TX_collision_detect_set => \TX_collision_detect_set\, 
        N_480_rs_0 => \N_480_rs_0\, un33_int_reg_clr => 
        un33_int_reg_clr, rx_CRC_error_set => \rx_CRC_error_set\, 
        N_480_rs => \N_480_rs\, un29_int_reg_clr => 
        un29_int_reg_clr, CommsFPGA_CCC_0_LOCK => 
        CommsFPGA_CCC_0_LOCK, CommsFPGA_top_0_INT => 
        CommsFPGA_top_0_INT, empty_r_3 => empty_r_3, N_357 => 
        N_357, tx_packet_complt => tx_packet_complt, DRVR_EN_c
         => \DRVR_EN_c\, N_209_i => N_209_i, rdiff_bus_cry_0_Y_0
         => rdiff_bus_cry_0_Y_0, N_314_i_i => N_314_i_i, m34 => 
        m34, un2_re_p_0 => un2_re_p, TX_FIFO_rd_en => 
        TX_FIFO_rd_en, CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, iRX_FIFO_rd_en_RNIJFNA_0
         => iRX_FIFO_rd_en_RNIJFNA_0, REN_d1_0 => REN_d1, N_283_i
         => N_283_i, N_6_0 => N_6_0, N_480 => N_480, 
        TX_PostAmble_d1 => TX_PostAmble_d1, RX_FIFO_RST_1 => 
        RX_FIFO_RST_1, RX_EarlyTerm => RX_EarlyTerm, 
        CoreAPB3_0_APBmslave0_PSELx => 
        CoreAPB3_0_APBmslave0_PSELx, un2_re_p => un2_re_p_0, 
        RX_FIFO_Empty => RX_FIFO_Empty, TX_FIFO_Full => 
        TX_FIFO_Full, RE_d1 => RE_d1, re_pulse_d1 => re_pulse_d1, 
        un19_tx_dataen => un19_tx_dataen, tx_preamble_pat_en => 
        tx_preamble_pat_en, TX_PreAmble => TX_PreAmble, 
        MANCHESTER_OUT_5 => MANCHESTER_OUT_5, BIT_CLK => 
        \BIT_CLK\, fifo_MEMRE => fifo_MEMRE, m35 => m35, 
        byte_clk_en => \byte_clk_en\, REN_d1 => REN_d1_0, 
        TX_FIFO_Empty => TX_FIFO_Empty, iTX_FIFO_rd_en => 
        iTX_FIFO_rd_en, RX_FIFO_Full => RX_FIFO_Full, 
        rx_packet_complt => rx_packet_complt, N_386_i_set => 
        \N_386_i_set\, un25_read_reg_en => un25_read_reg_en, 
        N_386_i_rs => \N_386_i_rs\, TX_FIFO_wr_en => 
        TX_FIFO_wr_en, N_209_i_i => N_209_i_i, RX_FIFO_rd_en => 
        RX_FIFO_rd_en, TX_FIFO_RST => TX_FIFO_RST, start_tx_FIFO
         => start_tx_FIFO, internal_loopback => internal_loopback, 
        long_reset => \long_reset\, CoreAPB3_0_APBmslave0_PREADY
         => CoreAPB3_0_APBmslave0_PREADY, long_reset_set => 
        \long_reset_set\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, long_reset_i => long_reset_i, 
        un2_apb3_addr_13 => un2_apb3_addr_13, N_386_i_i => 
        N_386_i_i, N_106_mux_i_i => N_106_mux_i_i);
    
    bd_reset_RNIK1J6 : CLKINT
      port map(A => \bd_reset\, Y => bd_reset_i);
    
    RX_FIFO_UNDERRUN_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un21_int_reg_clr, ALn => RX_FIFO_UNDERRUN_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_UNDERRUN_set\);
    
    \long_reset_cntr[4]\ : SLE
      port map(D => \long_reset_cntr_3[4]_net_1\, CLK => 
        \BIT_CLK\, EN => VCC_net_1, ALn => bd_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[4]_net_1\);
    
    N_386_i_rs : SLE
      port map(D => VCC_net_1, CLK => un2_apb3_addr_13, EN => 
        VCC_net_1, ALn => N_386_i_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \N_386_i_rs\);
    
    \ClkDivider[1]\ : SLE
      port map(D => \ClkDivider_RNO[1]_net_1\, CLK => \BIT_CLK\, 
        EN => VCC_net_1, ALn => bd_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ClkDivider[1]_net_1\);
    
    TX_collision_detect_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un33_int_reg_clr, ALn => TX_collision_detect_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \TX_collision_detect_set\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som is

    port( DEBOUNCE_IN           : in    std_logic_vector(2 downto 0);
          ID_RES                : in    std_logic_vector(3 downto 0);
          MAC_MII_RXD           : in    std_logic_vector(3 downto 0);
          MAC_MII_TXD           : out   std_logic_vector(3 downto 0);
          MDDR_ADDR             : out   std_logic_vector(15 downto 0);
          MDDR_BA               : out   std_logic_vector(2 downto 0);
          GPIO_1_BI             : inout std_logic_vector(0 to 0) := (others => 'Z');
          GPIO_1_BIDI           : in    std_logic_vector(0 to 0);
          GPIO_6_PAD            : inout std_logic_vector(0 to 0) := (others => 'Z');
          GPIO_7_PADI           : inout std_logic_vector(0 to 0) := (others => 'Z');
          MDDR_DM_RDQS          : inout std_logic_vector(1 downto 0) := (others => 'Z');
          MDDR_DQ               : inout std_logic_vector(15 downto 0) := (others => 'Z');
          MDDR_DQS              : inout std_logic_vector(1 downto 0) := (others => 'Z');
          SPI_1_CLK             : inout std_logic_vector(0 to 0) := (others => 'Z');
          SPI_1_SS0_CAM         : inout std_logic_vector(0 to 0) := (others => 'Z');
          SPI_1_SS0_OTH         : inout std_logic_vector(0 to 0) := (others => 'Z');
          DEVRST_N              : in    std_logic;
          MAC_MII_COL           : in    std_logic;
          MAC_MII_CRS           : in    std_logic;
          MAC_MII_RX_CLK        : in    std_logic;
          MAC_MII_RX_DV         : in    std_logic;
          MAC_MII_RX_ER         : in    std_logic;
          MAC_MII_TX_CLK        : in    std_logic;
          MANCHESTER_IN         : in    std_logic;
          MDDR_DQS_TMATCH_0_IN  : in    std_logic;
          MMUART_0_RXD_F2M      : in    std_logic;
          MMUART_1_RXD          : in    std_logic;
          PULLDOWN_R9           : in    std_logic;
          SPI_0_DI              : in    std_logic;
          SPI_1_DI_CAM          : in    std_logic;
          SPI_1_DI_OTH          : in    std_logic;
          XTL                   : in    std_logic;
          DEBOUNCE_OUT_1        : out   std_logic;
          DEBOUNCE_OUT_2        : out   std_logic;
          DRVR_EN               : out   std_logic;
          Data_FAIL             : out   std_logic;
          GPIO_11_M2F           : out   std_logic;
          GPIO_20_OUT           : out   std_logic;
          GPIO_21_M2F           : out   std_logic;
          GPIO_22_M2F           : out   std_logic;
          GPIO_24_M2F           : out   std_logic;
          GPIO_5_M2F            : out   std_logic;
          GPIO_8_M2F            : out   std_logic;
          MAC_MII_MDC           : out   std_logic;
          MAC_MII_TX_EN         : out   std_logic;
          MANCH_OUT_N           : out   std_logic;
          MANCH_OUT_P           : out   std_logic;
          MDDR_CAS_N            : out   std_logic;
          MDDR_CKE              : out   std_logic;
          MDDR_CLK              : out   std_logic;
          MDDR_CLK_N            : out   std_logic;
          MDDR_CS_N             : out   std_logic;
          MDDR_DQS_TMATCH_0_OUT : out   std_logic;
          MDDR_ODT              : out   std_logic;
          MDDR_RAS_N            : out   std_logic;
          MDDR_RESET_N          : out   std_logic;
          MDDR_WE_N             : out   std_logic;
          MMUART_0_TXD_M2F      : out   std_logic;
          MMUART_1_TXD          : out   std_logic;
          RCVR_EN               : out   std_logic;
          SPI_0_DO              : out   std_logic;
          SPI_0_SS1             : out   std_logic;
          SPI_1_DO_CAM          : out   std_logic;
          SPI_1_DO_OTH          : out   std_logic;
          GPIO_0_BI             : inout std_logic := 'Z';
          GPIO_12_BI            : inout std_logic := 'Z';
          GPIO_14_BI            : inout std_logic := 'Z';
          GPIO_15_BI            : inout std_logic := 'Z';
          GPIO_16_BI            : inout std_logic := 'Z';
          GPIO_17_BI            : inout std_logic := 'Z';
          GPIO_18_BI            : inout std_logic := 'Z';
          GPIO_25_BI            : inout std_logic := 'Z';
          GPIO_26_BI            : inout std_logic := 'Z';
          GPIO_31_BI            : inout std_logic := 'Z';
          GPIO_3_BI             : inout std_logic := 'Z';
          GPIO_4_BI             : inout std_logic := 'Z';
          I2C_1_SCL             : inout std_logic := 'Z';
          I2C_1_SDA             : inout std_logic := 'Z';
          MAC_MII_MDIO          : inout std_logic := 'Z';
          SPI_0_CLK             : inout std_logic := 'Z';
          SPI_0_SS0             : inout std_logic := 'Z'
        );

end m2s010_som;

architecture DEF_ARCH of m2s010_som is 

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component CoreAPB3
    port( m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(15 downto 12) := (others => 'U');
          CoreAPB3_0_APBmslave0_PSELx            : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component m2s010_som_CommsFPGA_CCC_0_FCCC
    port( m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : in    std_logic := 'U';
          CommsFPGA_CCC_0_LOCK                      : out   std_logic;
          CommsFPGA_CCC_0_GL1                       : out   std_logic;
          CommsFPGA_CCC_0_GL0                       : out   std_logic
        );
  end component;

  component m2s010_som_ID_RES_0_IO
    port( ID_RES  : in    std_logic_vector(3 downto 0) := (others => 'U');
          Y_net_0 : out   std_logic_vector(3 downto 0)
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component m2s010_som_sb
    port( MDDR_DQS                                  : inout   std_logic_vector(1 downto 0);
          MDDR_DQ                                   : inout   std_logic_vector(15 downto 0);
          MDDR_DM_RDQS                              : inout   std_logic_vector(1 downto 0);
          MDDR_BA                                   : out   std_logic_vector(2 downto 0);
          MDDR_ADDR                                 : out   std_logic_vector(15 downto 0);
          CoreAPB3_0_APBmslave0_PADDR               : out   std_logic_vector(7 downto 0);
          m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR    : out   std_logic_vector(15 downto 12);
          CoreAPB3_0_APBmslave0_PWDATA              : out   std_logic_vector(7 downto 0);
          MAC_MII_TXD_c                             : out   std_logic_vector(3 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA_m            : in    std_logic_vector(7 downto 0) := (others => 'U');
          Y_net_0                                   : in    std_logic_vector(3 downto 0) := (others => 'U');
          MAC_MII_RXD_c                             : in    std_logic_vector(3 downto 0) := (others => 'U');
          SPI_1_SS0_OTH_0                           : inout   std_logic;
          DEBOUNCE_OUT_net_0_0                      : in    std_logic := 'U';
          GPIO_7_PADI_0                             : inout   std_logic;
          GPIO_6_PAD_0                              : inout   std_logic;
          GPIO_1_BI_0                               : inout   std_logic;
          SPI_1_SS0_CAM_0                           : inout   std_logic;
          SPI_1_CLK_0                               : inout   std_logic;
          SPI_0_SS1                                 : out   std_logic;
          SPI_0_SS0                                 : inout   std_logic;
          SPI_0_DO                                  : out   std_logic;
          SPI_0_DI                                  : in    std_logic := 'U';
          SPI_0_CLK                                 : inout   std_logic;
          MMUART_1_TXD                              : out   std_logic;
          MMUART_1_RXD                              : in    std_logic := 'U';
          MDDR_WE_N                                 : out   std_logic;
          MDDR_RESET_N                              : out   std_logic;
          MDDR_RAS_N                                : out   std_logic;
          MDDR_ODT                                  : out   std_logic;
          MDDR_DQS_TMATCH_0_OUT                     : out   std_logic;
          MDDR_DQS_TMATCH_0_IN                      : in    std_logic := 'U';
          MDDR_CS_N                                 : out   std_logic;
          MDDR_CKE                                  : out   std_logic;
          MDDR_CAS_N                                : out   std_logic;
          I2C_1_SDA                                 : inout   std_logic;
          I2C_1_SCL                                 : inout   std_logic;
          GPIO_31_BI                                : inout   std_logic;
          GPIO_26_BI                                : inout   std_logic;
          GPIO_25_BI                                : inout   std_logic;
          GPIO_20_OUT                               : out   std_logic;
          GPIO_18_BI                                : inout   std_logic;
          GPIO_17_BI                                : inout   std_logic;
          GPIO_16_BI                                : inout   std_logic;
          GPIO_15_BI                                : inout   std_logic;
          GPIO_14_BI                                : inout   std_logic;
          GPIO_12_BI                                : inout   std_logic;
          GPIO_4_BI                                 : inout   std_logic;
          GPIO_3_BI                                 : inout   std_logic;
          GPIO_0_BI                                 : inout   std_logic;
          CoreAPB3_0_APBmslave0_PENABLE             : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx    : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE              : out   std_logic;
          MAC_MII_MDC_c                             : out   std_logic;
          GPIO_22_M2F_c                             : out   std_logic;
          GPIO_21_M2F_c                             : out   std_logic;
          m2s010_som_sb_0_GPIO_28_SW_RESET          : out   std_logic;
          MMUART_0_TXD_M2F_c                        : out   std_logic;
          GPIO_24_M2F_c                             : out   std_logic;
          GPIO_5_M2F_c                              : out   std_logic;
          GPIO_8_M2F_c                              : out   std_logic;
          GPIO_11_M2F_c                             : out   std_logic;
          MAC_MII_TX_EN_c                           : out   std_logic;
          MAC_MII_COL_c                             : in    std_logic := 'U';
          MAC_MII_CRS_c                             : in    std_logic := 'U';
          CommsFPGA_top_0_INT                       : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY_i_m_i        : in    std_logic := 'U';
          DEBOUNCE_OUT_1_c                          : in    std_logic := 'U';
          DEBOUNCE_OUT_2_c                          : in    std_logic := 'U';
          MMUART_0_RXD_F2M_c                        : in    std_logic := 'U';
          MAC_MII_RX_CLK_c                          : in    std_logic := 'U';
          MAC_MII_RX_DV_c                           : in    std_logic := 'U';
          MAC_MII_RX_ER_c                           : in    std_logic := 'U';
          MAC_MII_TX_CLK_c                          : in    std_logic := 'U';
          MDDR_CLK_N                                : out   std_logic;
          MDDR_CLK                                  : out   std_logic;
          XTL                                       : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz                 : out   std_logic;
          m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : inout   std_logic;
          SPI_1_DI_CAM_c                            : in    std_logic := 'U';
          SPI_1_DI_OTH_c                            : in    std_logic := 'U';
          CommsFPGA_top_0_CAMERA_NODE               : in    std_logic := 'U';
          DEVRST_N                                  : in    std_logic := 'U';
          m2s010_som_sb_0_POWER_ON_RESET_N          : out   std_logic;
          MAC_MII_MDIO                              : inout   std_logic;
          SPI_1_DO_CAM_c                            : inout   std_logic;
          SPI_1_DO_OTH                              : out   std_logic
        );
  end component;

  component CommsFPGA_top
    port( CoreAPB3_0_APBmslave0_PWDATA       : in    std_logic_vector(7 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PRDATA_m     : out   std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PADDR        : in    std_logic_vector(7 downto 0) := (others => 'U');
          DEBOUNCE_IN_c                      : in    std_logic_vector(2 downto 0) := (others => 'U');
          Y_net_0                            : in    std_logic_vector(3 downto 1) := (others => 'U');
          DEBOUNCE_OUT_net_0_0               : out   std_logic;
          MANCHESTER_IN_c                    : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY_i_m_i : out   std_logic;
          MANCH_OUT_P_c                      : out   std_logic;
          MANCH_OUT_P_c_i                    : out   std_logic;
          N_209_i_i                          : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PSELx        : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PWRITE       : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PENABLE      : in    std_logic := 'U';
          N_209_i                            : out   std_logic;
          DRVR_EN_c                          : out   std_logic;
          CommsFPGA_top_0_INT                : out   std_logic;
          CommsFPGA_CCC_0_LOCK               : in    std_logic := 'U';
          DEBOUNCE_OUT_1_c                   : out   std_logic;
          DEBOUNCE_OUT_2_c                   : out   std_logic;
          CommsFPGA_top_0_CAMERA_NODE        : out   std_logic;
          m2s010_som_sb_0_POWER_ON_RESET_N   : in    std_logic := 'U';
          m2s010_som_sb_0_GPIO_28_SW_RESET   : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL1                : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0                : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz          : in    std_logic := 'U'
        );
  end component;

    signal m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC, 
        CommsFPGA_CCC_0_LOCK, CommsFPGA_CCC_0_GL0, 
        CommsFPGA_CCC_0_GL1, m2s010_som_sb_0_GPIO_28_SW_RESET, 
        m2s010_som_sb_0_POWER_ON_RESET_N, 
        m2s010_som_sb_0_CCC_71MHz, \Y_net_0[0]\, \Y_net_0[1]\, 
        \Y_net_0[2]\, \Y_net_0[3]\, CommsFPGA_top_0_CAMERA_NODE, 
        CommsFPGA_top_0_INT, \DEBOUNCE_OUT_net_0[0]\, GND_net_1, 
        \CoreAPB3_0_APBmslave0_PADDR[0]\, 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, 
        \CoreAPB3_0_APBmslave0_PADDR[5]\, 
        \CoreAPB3_0_APBmslave0_PADDR[6]\, 
        \CoreAPB3_0_APBmslave0_PADDR[7]\, 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[12]\, 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[13]\, 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[14]\, 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[15]\, 
        CoreAPB3_0_APBmslave0_PWRITE, 
        CoreAPB3_0_APBmslave0_PENABLE, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx, 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, VCC_net_1, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[0]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[1]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[2]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[3]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[4]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[5]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[6]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[7]\, 
        CoreAPB3_0_APBmslave0_PSELx, \DEBOUNCE_IN_c[0]\, 
        \DEBOUNCE_IN_c[1]\, \DEBOUNCE_IN_c[2]\, MAC_MII_COL_c, 
        MAC_MII_CRS_c, \MAC_MII_RXD_c[0]\, \MAC_MII_RXD_c[1]\, 
        \MAC_MII_RXD_c[2]\, \MAC_MII_RXD_c[3]\, MAC_MII_RX_CLK_c, 
        MAC_MII_RX_DV_c, MAC_MII_RX_ER_c, MAC_MII_TX_CLK_c, 
        MANCHESTER_IN_c, MMUART_0_RXD_F2M_c, Data_FAIL_c, 
        SPI_1_DI_CAM_c, SPI_1_DI_OTH_c, DEBOUNCE_OUT_1_c, 
        DEBOUNCE_OUT_2_c, DRVR_EN_c, GPIO_11_M2F_c, GPIO_21_M2F_c, 
        GPIO_22_M2F_c, GPIO_24_M2F_c, GPIO_5_M2F_c, GPIO_8_M2F_c, 
        MAC_MII_MDC_c, \MAC_MII_TXD_c[0]\, \MAC_MII_TXD_c[1]\, 
        \MAC_MII_TXD_c[2]\, \MAC_MII_TXD_c[3]\, MAC_MII_TX_EN_c, 
        MANCH_OUT_P_c, MMUART_0_TXD_M2F_c, SPI_1_DO_CAM_c, 
        MANCH_OUT_P_c_i, CoreAPB3_0_APBmslave0_PREADY_i_m_i, 
        \CommsFPGA_top_0.N_209_i_i\, N_209_i : std_logic;

    for all : CoreAPB3
	Use entity work.CoreAPB3(DEF_ARCH);
    for all : m2s010_som_CommsFPGA_CCC_0_FCCC
	Use entity work.m2s010_som_CommsFPGA_CCC_0_FCCC(DEF_ARCH);
    for all : m2s010_som_ID_RES_0_IO
	Use entity work.m2s010_som_ID_RES_0_IO(DEF_ARCH);
    for all : m2s010_som_sb
	Use entity work.m2s010_som_sb(DEF_ARCH);
    for all : CommsFPGA_top
	Use entity work.CommsFPGA_top(DEF_ARCH);
begin 


    RCVR_EN_obuf : OUTBUF
      port map(D => VCC_net_1, PAD => RCVR_EN);
    
    MANCH_OUT_N_obuf : OUTBUF
      port map(D => MANCH_OUT_P_c_i, PAD => MANCH_OUT_N);
    
    \MAC_MII_RXD_ibuf[1]\ : INBUF
      port map(PAD => MAC_MII_RXD(1), Y => \MAC_MII_RXD_c[1]\);
    
    MMUART_0_RXD_F2M_ibuf : INBUF
      port map(PAD => MMUART_0_RXD_F2M, Y => MMUART_0_RXD_F2M_c);
    
    MAC_MII_RX_CLK_ibuf : INBUF
      port map(PAD => MAC_MII_RX_CLK, Y => MAC_MII_RX_CLK_c);
    
    MAC_MII_CRS_ibuf : INBUF
      port map(PAD => MAC_MII_CRS, Y => MAC_MII_CRS_c);
    
    CoreAPB3_0 : CoreAPB3
      port map(m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[15]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[14]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[13]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[12]\, 
        CoreAPB3_0_APBmslave0_PSELx => 
        CoreAPB3_0_APBmslave0_PSELx, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    CommsFPGA_CCC_0 : m2s010_som_CommsFPGA_CCC_0_FCCC
      port map(m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC, 
        CommsFPGA_CCC_0_LOCK => CommsFPGA_CCC_0_LOCK, 
        CommsFPGA_CCC_0_GL1 => CommsFPGA_CCC_0_GL1, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0);
    
    MAC_MII_TX_EN_obuf : OUTBUF
      port map(D => MAC_MII_TX_EN_c, PAD => MAC_MII_TX_EN);
    
    MAC_MII_TX_CLK_ibuf : INBUF
      port map(PAD => MAC_MII_TX_CLK, Y => MAC_MII_TX_CLK_c);
    
    \MAC_MII_TXD_obuf[1]\ : OUTBUF
      port map(D => \MAC_MII_TXD_c[1]\, PAD => MAC_MII_TXD(1));
    
    DEBOUNCE_OUT_2_obuf : OUTBUF
      port map(D => DEBOUNCE_OUT_2_c, PAD => DEBOUNCE_OUT_2);
    
    ID_RES_0 : m2s010_som_ID_RES_0_IO
      port map(ID_RES(3) => ID_RES(3), ID_RES(2) => ID_RES(2), 
        ID_RES(1) => ID_RES(1), ID_RES(0) => ID_RES(0), 
        Y_net_0(3) => \Y_net_0[3]\, Y_net_0(2) => \Y_net_0[2]\, 
        Y_net_0(1) => \Y_net_0[1]\, Y_net_0(0) => \Y_net_0[0]\);
    
    \MAC_MII_RXD_ibuf[0]\ : INBUF
      port map(PAD => MAC_MII_RXD(0), Y => \MAC_MII_RXD_c[0]\);
    
    MMUART_0_TXD_M2F_obuf : OUTBUF
      port map(D => MMUART_0_TXD_M2F_c, PAD => MMUART_0_TXD_M2F);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \MAC_MII_RXD_ibuf[3]\ : INBUF
      port map(PAD => MAC_MII_RXD(3), Y => \MAC_MII_RXD_c[3]\);
    
    SPI_1_DI_CAM_ibuf : INBUF
      port map(PAD => SPI_1_DI_CAM, Y => SPI_1_DI_CAM_c);
    
    \MAC_MII_TXD_obuf[0]\ : OUTBUF
      port map(D => \MAC_MII_TXD_c[0]\, PAD => MAC_MII_TXD(0));
    
    Data_FAIL_obuf : OUTBUF
      port map(D => Data_FAIL_c, PAD => Data_FAIL);
    
    MAC_MII_COL_ibuf : INBUF
      port map(PAD => MAC_MII_COL, Y => MAC_MII_COL_c);
    
    I_291 : CLKINT
      port map(A => N_209_i, Y => \CommsFPGA_top_0.N_209_i_i\);
    
    MANCH_OUT_P_obuf : OUTBUF
      port map(D => MANCH_OUT_P_c, PAD => MANCH_OUT_P);
    
    MAC_MII_MDC_obuf : OUTBUF
      port map(D => MAC_MII_MDC_c, PAD => MAC_MII_MDC);
    
    MANCHESTER_IN_ibuf : INBUF
      port map(PAD => MANCHESTER_IN, Y => MANCHESTER_IN_c);
    
    GPIO_22_M2F_obuf : OUTBUF
      port map(D => GPIO_22_M2F_c, PAD => GPIO_22_M2F);
    
    GPIO_21_M2F_obuf : OUTBUF
      port map(D => GPIO_21_M2F_c, PAD => GPIO_21_M2F);
    
    SPI_1_DO_CAM_obuf : OUTBUF
      port map(D => SPI_1_DO_CAM_c, PAD => SPI_1_DO_CAM);
    
    \MAC_MII_TXD_obuf[3]\ : OUTBUF
      port map(D => \MAC_MII_TXD_c[3]\, PAD => MAC_MII_TXD(3));
    
    \DEBOUNCE_IN_ibuf[1]\ : INBUF
      port map(PAD => DEBOUNCE_IN(1), Y => \DEBOUNCE_IN_c[1]\);
    
    MAC_MII_RX_DV_ibuf : INBUF
      port map(PAD => MAC_MII_RX_DV, Y => MAC_MII_RX_DV_c);
    
    DRVR_EN_obuf : OUTBUF
      port map(D => DRVR_EN_c, PAD => DRVR_EN);
    
    DEBOUNCE_OUT_1_obuf : OUTBUF
      port map(D => DEBOUNCE_OUT_1_c, PAD => DEBOUNCE_OUT_1);
    
    SPI_1_DI_OTH_ibuf : INBUF
      port map(PAD => SPI_1_DI_OTH, Y => SPI_1_DI_OTH_c);
    
    m2s010_som_sb_0 : m2s010_som_sb
      port map(MDDR_DQS(1) => MDDR_DQS(1), MDDR_DQS(0) => 
        MDDR_DQS(0), MDDR_DQ(15) => MDDR_DQ(15), MDDR_DQ(14) => 
        MDDR_DQ(14), MDDR_DQ(13) => MDDR_DQ(13), MDDR_DQ(12) => 
        MDDR_DQ(12), MDDR_DQ(11) => MDDR_DQ(11), MDDR_DQ(10) => 
        MDDR_DQ(10), MDDR_DQ(9) => MDDR_DQ(9), MDDR_DQ(8) => 
        MDDR_DQ(8), MDDR_DQ(7) => MDDR_DQ(7), MDDR_DQ(6) => 
        MDDR_DQ(6), MDDR_DQ(5) => MDDR_DQ(5), MDDR_DQ(4) => 
        MDDR_DQ(4), MDDR_DQ(3) => MDDR_DQ(3), MDDR_DQ(2) => 
        MDDR_DQ(2), MDDR_DQ(1) => MDDR_DQ(1), MDDR_DQ(0) => 
        MDDR_DQ(0), MDDR_DM_RDQS(1) => MDDR_DM_RDQS(1), 
        MDDR_DM_RDQS(0) => MDDR_DM_RDQS(0), MDDR_BA(2) => 
        MDDR_BA(2), MDDR_BA(1) => MDDR_BA(1), MDDR_BA(0) => 
        MDDR_BA(0), MDDR_ADDR(15) => MDDR_ADDR(15), MDDR_ADDR(14)
         => MDDR_ADDR(14), MDDR_ADDR(13) => MDDR_ADDR(13), 
        MDDR_ADDR(12) => MDDR_ADDR(12), MDDR_ADDR(11) => 
        MDDR_ADDR(11), MDDR_ADDR(10) => MDDR_ADDR(10), 
        MDDR_ADDR(9) => MDDR_ADDR(9), MDDR_ADDR(8) => 
        MDDR_ADDR(8), MDDR_ADDR(7) => MDDR_ADDR(7), MDDR_ADDR(6)
         => MDDR_ADDR(6), MDDR_ADDR(5) => MDDR_ADDR(5), 
        MDDR_ADDR(4) => MDDR_ADDR(4), MDDR_ADDR(3) => 
        MDDR_ADDR(3), MDDR_ADDR(2) => MDDR_ADDR(2), MDDR_ADDR(1)
         => MDDR_ADDR(1), MDDR_ADDR(0) => MDDR_ADDR(0), 
        CoreAPB3_0_APBmslave0_PADDR(7) => 
        \CoreAPB3_0_APBmslave0_PADDR[7]\, 
        CoreAPB3_0_APBmslave0_PADDR(6) => 
        \CoreAPB3_0_APBmslave0_PADDR[6]\, 
        CoreAPB3_0_APBmslave0_PADDR(5) => 
        \CoreAPB3_0_APBmslave0_PADDR[5]\, 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        \CoreAPB3_0_APBmslave0_PADDR[0]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[15]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[14]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[13]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[12]\, 
        CoreAPB3_0_APBmslave0_PWDATA(7) => 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, MAC_MII_TXD_c(3) => 
        \MAC_MII_TXD_c[3]\, MAC_MII_TXD_c(2) => 
        \MAC_MII_TXD_c[2]\, MAC_MII_TXD_c(1) => 
        \MAC_MII_TXD_c[1]\, MAC_MII_TXD_c(0) => 
        \MAC_MII_TXD_c[0]\, CoreAPB3_0_APBmslave0_PRDATA_m(7) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[7]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(6) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[6]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(5) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[5]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(4) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[4]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(3) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[3]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(2) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[2]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(1) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[1]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(0) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[0]\, Y_net_0(3) => 
        \Y_net_0[3]\, Y_net_0(2) => \Y_net_0[2]\, Y_net_0(1) => 
        \Y_net_0[1]\, Y_net_0(0) => \Y_net_0[0]\, 
        MAC_MII_RXD_c(3) => \MAC_MII_RXD_c[3]\, MAC_MII_RXD_c(2)
         => \MAC_MII_RXD_c[2]\, MAC_MII_RXD_c(1) => 
        \MAC_MII_RXD_c[1]\, MAC_MII_RXD_c(0) => 
        \MAC_MII_RXD_c[0]\, SPI_1_SS0_OTH_0 => SPI_1_SS0_OTH(0), 
        DEBOUNCE_OUT_net_0_0 => \DEBOUNCE_OUT_net_0[0]\, 
        GPIO_7_PADI_0 => GPIO_7_PADI(0), GPIO_6_PAD_0 => 
        GPIO_6_PAD(0), GPIO_1_BI_0 => GPIO_1_BI(0), 
        SPI_1_SS0_CAM_0 => SPI_1_SS0_CAM(0), SPI_1_CLK_0 => 
        SPI_1_CLK(0), SPI_0_SS1 => SPI_0_SS1, SPI_0_SS0 => 
        SPI_0_SS0, SPI_0_DO => SPI_0_DO, SPI_0_DI => SPI_0_DI, 
        SPI_0_CLK => SPI_0_CLK, MMUART_1_TXD => MMUART_1_TXD, 
        MMUART_1_RXD => MMUART_1_RXD, MDDR_WE_N => MDDR_WE_N, 
        MDDR_RESET_N => MDDR_RESET_N, MDDR_RAS_N => MDDR_RAS_N, 
        MDDR_ODT => MDDR_ODT, MDDR_DQS_TMATCH_0_OUT => 
        MDDR_DQS_TMATCH_0_OUT, MDDR_DQS_TMATCH_0_IN => 
        MDDR_DQS_TMATCH_0_IN, MDDR_CS_N => MDDR_CS_N, MDDR_CKE
         => MDDR_CKE, MDDR_CAS_N => MDDR_CAS_N, I2C_1_SDA => 
        I2C_1_SDA, I2C_1_SCL => I2C_1_SCL, GPIO_31_BI => 
        GPIO_31_BI, GPIO_26_BI => GPIO_26_BI, GPIO_25_BI => 
        GPIO_25_BI, GPIO_20_OUT => GPIO_20_OUT, GPIO_18_BI => 
        GPIO_18_BI, GPIO_17_BI => GPIO_17_BI, GPIO_16_BI => 
        GPIO_16_BI, GPIO_15_BI => GPIO_15_BI, GPIO_14_BI => 
        GPIO_14_BI, GPIO_12_BI => GPIO_12_BI, GPIO_4_BI => 
        GPIO_4_BI, GPIO_3_BI => GPIO_3_BI, GPIO_0_BI => GPIO_0_BI, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, MAC_MII_MDC_c => 
        MAC_MII_MDC_c, GPIO_22_M2F_c => GPIO_22_M2F_c, 
        GPIO_21_M2F_c => GPIO_21_M2F_c, 
        m2s010_som_sb_0_GPIO_28_SW_RESET => 
        m2s010_som_sb_0_GPIO_28_SW_RESET, MMUART_0_TXD_M2F_c => 
        MMUART_0_TXD_M2F_c, GPIO_24_M2F_c => GPIO_24_M2F_c, 
        GPIO_5_M2F_c => GPIO_5_M2F_c, GPIO_8_M2F_c => 
        GPIO_8_M2F_c, GPIO_11_M2F_c => GPIO_11_M2F_c, 
        MAC_MII_TX_EN_c => MAC_MII_TX_EN_c, MAC_MII_COL_c => 
        MAC_MII_COL_c, MAC_MII_CRS_c => MAC_MII_CRS_c, 
        CommsFPGA_top_0_INT => CommsFPGA_top_0_INT, 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, DEBOUNCE_OUT_1_c => 
        DEBOUNCE_OUT_1_c, DEBOUNCE_OUT_2_c => DEBOUNCE_OUT_2_c, 
        MMUART_0_RXD_F2M_c => MMUART_0_RXD_F2M_c, 
        MAC_MII_RX_CLK_c => MAC_MII_RX_CLK_c, MAC_MII_RX_DV_c => 
        MAC_MII_RX_DV_c, MAC_MII_RX_ER_c => MAC_MII_RX_ER_c, 
        MAC_MII_TX_CLK_c => MAC_MII_TX_CLK_c, MDDR_CLK_N => 
        MDDR_CLK_N, MDDR_CLK => MDDR_CLK, XTL => XTL, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC, SPI_1_DI_CAM_c
         => SPI_1_DI_CAM_c, SPI_1_DI_OTH_c => SPI_1_DI_OTH_c, 
        CommsFPGA_top_0_CAMERA_NODE => 
        CommsFPGA_top_0_CAMERA_NODE, DEVRST_N => DEVRST_N, 
        m2s010_som_sb_0_POWER_ON_RESET_N => 
        m2s010_som_sb_0_POWER_ON_RESET_N, MAC_MII_MDIO => 
        MAC_MII_MDIO, SPI_1_DO_CAM_c => SPI_1_DO_CAM_c, 
        SPI_1_DO_OTH => SPI_1_DO_OTH);
    
    GPIO_24_M2F_obuf : OUTBUF
      port map(D => GPIO_24_M2F_c, PAD => GPIO_24_M2F);
    
    \DEBOUNCE_IN_ibuf[2]\ : INBUF
      port map(PAD => DEBOUNCE_IN(2), Y => \DEBOUNCE_IN_c[2]\);
    
    \MAC_MII_RXD_ibuf[2]\ : INBUF
      port map(PAD => MAC_MII_RXD(2), Y => \MAC_MII_RXD_c[2]\);
    
    PULLDOWN_R9_ibuf : INBUF
      port map(PAD => PULLDOWN_R9, Y => Data_FAIL_c);
    
    GPIO_11_M2F_obuf : OUTBUF
      port map(D => GPIO_11_M2F_c, PAD => GPIO_11_M2F);
    
    GPIO_8_M2F_obuf : OUTBUF
      port map(D => GPIO_8_M2F_c, PAD => GPIO_8_M2F);
    
    \MAC_MII_TXD_obuf[2]\ : OUTBUF
      port map(D => \MAC_MII_TXD_c[2]\, PAD => MAC_MII_TXD(2));
    
    MAC_MII_RX_ER_ibuf : INBUF
      port map(PAD => MAC_MII_RX_ER, Y => MAC_MII_RX_ER_c);
    
    \DEBOUNCE_IN_ibuf[0]\ : INBUF
      port map(PAD => DEBOUNCE_IN(0), Y => \DEBOUNCE_IN_c[0]\);
    
    GPIO_5_M2F_obuf : OUTBUF
      port map(D => GPIO_5_M2F_c, PAD => GPIO_5_M2F);
    
    CommsFPGA_top_0 : CommsFPGA_top
      port map(CoreAPB3_0_APBmslave0_PWDATA(7) => 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(7) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[7]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(6) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[6]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(5) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[5]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(4) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[4]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(3) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[3]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(2) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[2]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(1) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[1]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(0) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[0]\, 
        CoreAPB3_0_APBmslave0_PADDR(7) => 
        \CoreAPB3_0_APBmslave0_PADDR[7]\, 
        CoreAPB3_0_APBmslave0_PADDR(6) => 
        \CoreAPB3_0_APBmslave0_PADDR[6]\, 
        CoreAPB3_0_APBmslave0_PADDR(5) => 
        \CoreAPB3_0_APBmslave0_PADDR[5]\, 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        \CoreAPB3_0_APBmslave0_PADDR[0]\, DEBOUNCE_IN_c(2) => 
        \DEBOUNCE_IN_c[2]\, DEBOUNCE_IN_c(1) => 
        \DEBOUNCE_IN_c[1]\, DEBOUNCE_IN_c(0) => 
        \DEBOUNCE_IN_c[0]\, Y_net_0(3) => \Y_net_0[3]\, 
        Y_net_0(2) => \Y_net_0[2]\, Y_net_0(1) => \Y_net_0[1]\, 
        DEBOUNCE_OUT_net_0_0 => \DEBOUNCE_OUT_net_0[0]\, 
        MANCHESTER_IN_c => MANCHESTER_IN_c, 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, MANCH_OUT_P_c => 
        MANCH_OUT_P_c, MANCH_OUT_P_c_i => MANCH_OUT_P_c_i, 
        N_209_i_i => \CommsFPGA_top_0.N_209_i_i\, 
        CoreAPB3_0_APBmslave0_PSELx => 
        CoreAPB3_0_APBmslave0_PSELx, CoreAPB3_0_APBmslave0_PWRITE
         => CoreAPB3_0_APBmslave0_PWRITE, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, N_209_i => N_209_i, 
        DRVR_EN_c => DRVR_EN_c, CommsFPGA_top_0_INT => 
        CommsFPGA_top_0_INT, CommsFPGA_CCC_0_LOCK => 
        CommsFPGA_CCC_0_LOCK, DEBOUNCE_OUT_1_c => 
        DEBOUNCE_OUT_1_c, DEBOUNCE_OUT_2_c => DEBOUNCE_OUT_2_c, 
        CommsFPGA_top_0_CAMERA_NODE => 
        CommsFPGA_top_0_CAMERA_NODE, 
        m2s010_som_sb_0_POWER_ON_RESET_N => 
        m2s010_som_sb_0_POWER_ON_RESET_N, 
        m2s010_som_sb_0_GPIO_28_SW_RESET => 
        m2s010_som_sb_0_GPIO_28_SW_RESET, CommsFPGA_CCC_0_GL1 => 
        CommsFPGA_CCC_0_GL1, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz);
    

end DEF_ARCH; 
